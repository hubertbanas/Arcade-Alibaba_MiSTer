library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity GFX1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of GFX1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"33",X"33",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"77",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"77",X"77",X"77",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"77",X"66",X"66",X"66",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"33",X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"11",X"33",X"33",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"77",X"77",X"77",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"33",X"33",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"77",X"77",X"77",X"77",X"77",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"00",X"00",X"08",X"0C",X"0C",X"08",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"01",X"00",X"00",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"0C",X"0E",X"0F",X"0F",X"0F",X"0F",X"0E",X"0C",X"03",X"07",X"0F",X"0F",X"0F",X"0F",X"07",X"03",
		X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"88",X"88",X"CC",X"EE",X"FF",X"FF",X"77",X"11",
		X"FF",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"EE",X"CC",X"88",X"88",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"11",X"77",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"66",X"66",X"66",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"33",X"BB",X"FF",X"EE",X"66",X"66",X"66",X"66",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"33",X"77",X"11",X"00",X"00",X"00",X"00",X"00",X"EE",
		X"11",X"11",X"11",X"11",X"11",X"11",X"FF",X"FF",X"00",X"00",X"88",X"88",X"CC",X"EE",X"FF",X"FF",
		X"00",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"33",
		X"EE",X"CC",X"CC",X"88",X"88",X"00",X"00",X"00",X"33",X"33",X"33",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",
		X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"77",X"77",X"33",X"22",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"DD",X"00",X"EE",X"DD",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",
		X"66",X"66",X"66",X"66",X"66",X"66",X"66",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"11",X"33",X"33",X"BB",X"FF",X"EE",X"00",X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"00",
		X"11",X"11",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"CC",X"EE",X"FF",X"FF",X"77",X"11",X"00",X"00",
		X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"CC",X"88",X"88",X"00",X"00",X"00",X"88",X"88",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"11",X"00",X"00",X"00",X"11",X"77",X"FF",X"FF",X"EE",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"88",X"88",X"88",X"88",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"CC",X"22",X"22",X"66",X"CC",X"88",X"00",X"33",X"77",X"CC",X"88",X"88",X"77",X"33",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"FF",X"FF",X"44",X"00",X"00",X"00",
		X"22",X"22",X"AA",X"AA",X"EE",X"EE",X"66",X"00",X"66",X"FF",X"BB",X"99",X"99",X"CC",X"44",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"88",X"DD",X"FF",X"BB",X"99",X"88",X"00",X"00",
		X"88",X"EE",X"EE",X"88",X"88",X"88",X"88",X"00",X"00",X"FF",X"FF",X"CC",X"66",X"33",X"11",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"11",X"BB",X"AA",X"AA",X"AA",X"EE",X"EE",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"00",X"99",X"99",X"99",X"DD",X"77",X"33",X"00",
		X"00",X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"CC",X"EE",X"BB",X"99",X"88",X"CC",X"CC",X"00",
		X"CC",X"EE",X"AA",X"AA",X"22",X"22",X"CC",X"00",X"00",X"66",X"99",X"99",X"BB",X"FF",X"66",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"22",X"00",X"00",X"77",X"FF",X"99",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"00",X"00",X"88",X"44",X"22",X"00",X"88",X"44",X"22",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",
		X"FF",X"77",X"33",X"33",X"33",X"33",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"33",X"33",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"88",X"88",X"88",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"CC",X"77",X"33",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"EE",X"00",X"66",X"FF",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"44",X"66",X"22",X"22",X"66",X"CC",X"88",X"00",X"44",X"CC",X"88",X"88",X"CC",X"77",X"33",X"00",
		X"88",X"CC",X"66",X"22",X"22",X"EE",X"EE",X"00",X"33",X"77",X"CC",X"88",X"88",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"88",X"99",X"99",X"99",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"00",X"88",X"99",X"99",X"99",X"99",X"FF",X"FF",X"00",
		X"EE",X"EE",X"22",X"22",X"66",X"CC",X"88",X"00",X"99",X"99",X"99",X"88",X"CC",X"77",X"33",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"11",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"EE",X"EE",X"22",X"22",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"88",X"CC",X"66",X"33",X"11",X"FF",X"FF",X"00",
		X"22",X"22",X"22",X"22",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",
		X"EE",X"EE",X"00",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"77",X"33",X"77",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"00",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"77",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"00",X"88",X"88",X"88",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"FF",X"00",
		X"AA",X"CC",X"EE",X"AA",X"22",X"EE",X"CC",X"00",X"77",X"FF",X"88",X"88",X"88",X"FF",X"77",X"00",
		X"22",X"66",X"EE",X"CC",X"88",X"EE",X"EE",X"00",X"77",X"FF",X"99",X"88",X"88",X"FF",X"FF",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"66",X"44",X"00",X"00",X"55",X"DD",X"99",X"99",X"FF",X"66",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"88",X"88",X"FF",X"FF",X"88",X"88",X"00",X"00",
		X"CC",X"EE",X"22",X"22",X"22",X"EE",X"CC",X"00",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"00",
		X"00",X"88",X"CC",X"EE",X"CC",X"88",X"00",X"00",X"FF",X"FF",X"11",X"00",X"11",X"FF",X"FF",X"00",
		X"EE",X"EE",X"CC",X"88",X"CC",X"EE",X"EE",X"00",X"FF",X"FF",X"11",X"33",X"11",X"FF",X"FF",X"00",
		X"66",X"EE",X"CC",X"88",X"CC",X"EE",X"66",X"00",X"CC",X"EE",X"77",X"33",X"77",X"EE",X"CC",X"00",
		X"00",X"00",X"EE",X"EE",X"00",X"00",X"00",X"00",X"EE",X"FF",X"11",X"11",X"FF",X"EE",X"00",X"00",
		X"22",X"22",X"22",X"AA",X"EE",X"EE",X"66",X"00",X"CC",X"EE",X"FF",X"BB",X"99",X"88",X"88",X"00",
		X"00",X"00",X"00",X"00",X"88",X"22",X"00",X"00",X"00",X"CC",X"EE",X"FF",X"33",X"00",X"00",X"00",
		X"CC",X"22",X"11",X"55",X"55",X"99",X"22",X"CC",X"33",X"44",X"88",X"AA",X"AA",X"99",X"44",X"33",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"EE",X"22",X"22",X"00",X"11",X"22",X"22",X"22",X"33",
		X"AA",X"AA",X"AA",X"22",X"00",X"00",X"00",X"EE",X"22",X"22",X"22",X"11",X"00",X"22",X"22",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"33",X"33",X"FF",X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",
		X"EE",X"EE",X"77",X"33",X"33",X"33",X"33",X"33",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"CC",X"CC",X"FF",X"FF",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",
		X"FF",X"FF",X"FF",X"33",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"CC",X"CC",X"EE",X"EE",X"77",X"33",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"88",X"88",X"FF",X"FF",X"FF",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"11",X"11",X"11",X"11",X"11",X"77",X"FF",X"FF",X"EE",X"CC",X"88",X"88",X"00",
		X"00",X"00",X"88",X"EE",X"EE",X"FF",X"FF",X"FF",X"00",X"00",X"11",X"77",X"77",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"88",X"88",X"88",X"DD",X"00",X"00",X"00",X"77",X"FF",X"DD",X"88",X"88",X"88",X"CC",X"66",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"CC",X"66",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"77",X"FF",X"DD",X"88",
		X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",
		X"CC",X"CC",X"CC",X"66",X"FF",X"FF",X"FF",X"CC",X"11",X"11",X"00",X"00",X"00",X"00",X"11",X"11",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",
		X"CC",X"CC",X"66",X"FF",X"FF",X"FF",X"00",X"EE",X"11",X"00",X"00",X"11",X"11",X"11",X"00",X"00",
		X"00",X"00",X"00",X"88",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"77",
		X"EE",X"EE",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"77",X"77",X"33",X"33",X"33",X"33",X"33",X"33",
		X"FF",X"FF",X"77",X"00",X"00",X"FF",X"FF",X"FF",X"11",X"00",X"00",X"00",X"00",X"11",X"11",X"11",
		X"88",X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"FF",X"FF",X"EE",X"00",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"22",X"CC",X"00",X"22",X"EE",X"22",X"00",X"00",X"88",X"77",X"00",X"00",X"FF",X"44",X"00",X"00",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"22",X"44",X"88",X"77",X"00",X"88",X"DD",X"AA",X"88",X"88",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"22",X"44",X"88",X"77",X"00",X"99",X"AA",X"AA",X"AA",X"EE",
		X"22",X"CC",X"00",X"00",X"00",X"EE",X"00",X"00",X"88",X"77",X"00",X"CC",X"BB",X"88",X"88",X"CC",
		X"00",X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"00",X"77",X"88",X"88",X"77",X"00",X"77",X"88",
		X"CC",X"22",X"22",X"CC",X"00",X"22",X"EE",X"22",X"77",X"88",X"88",X"77",X"00",X"00",X"FF",X"44",
		X"66",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"22",X"22",X"AA",X"77",X"88",X"88",X"77",X"00",X"66",X"99",X"88",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"88",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"77",X"88",X"88",X"77",X"00",X"88",X"DD",X"AA",
		X"22",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",
		X"CC",X"22",X"22",X"CC",X"00",X"CC",X"22",X"22",X"77",X"88",X"88",X"77",X"00",X"99",X"AA",X"AA",
		X"22",X"CC",X"00",X"CC",X"22",X"22",X"CC",X"00",X"88",X"77",X"00",X"77",X"88",X"88",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"88",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"07",X"0F",X"2D",X"2D",X"78",X"2D",X"00",X"00",X"00",X"04",X"06",X"06",X"07",X"07",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"2D",X"78",X"2D",X"3C",X"0F",X"07",X"03",X"00",X"07",X"07",X"06",X"06",X"04",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"04",X"06",X"06",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",X"00",X"03",X"07",X"0F",X"2D",X"2D",X"78",X"2D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"66",X"EE",X"6E",X"08",X"08",
		X"07",X"07",X"06",X"06",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"A5",X"F0",X"A5",X"A5",X"0F",X"3F",X"3F",X"00",X"2D",X"78",X"2D",X"3C",X"0F",X"07",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"08",X"4C",X"4C",X"44",X"EE",X"EE",X"00",
		X"00",X"77",X"FF",X"FF",X"9F",X"9F",X"FF",X"FF",X"00",X"30",X"70",X"70",X"70",X"F0",X"96",X"96",
		X"00",X"22",X"22",X"EE",X"EE",X"88",X"88",X"88",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",
		X"9F",X"9F",X"FF",X"FF",X"77",X"11",X"FF",X"00",X"F0",X"70",X"70",X"70",X"30",X"77",X"77",X"77",
		X"88",X"EE",X"EE",X"22",X"22",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",
		X"00",X"70",X"F0",X"F0",X"F0",X"F7",X"F7",X"F2",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"66",X"66",X"66",X"E6",X"E6",X"80",X"88",X"00",X"C0",X"E0",X"F0",X"87",X"A5",X"A5",X"B7",
		X"F2",X"F7",X"F7",X"F0",X"F0",X"F0",X"70",X"00",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",
		X"88",X"80",X"E6",X"E6",X"66",X"66",X"66",X"00",X"B7",X"A5",X"A5",X"87",X"F0",X"E0",X"C0",X"00",
		X"00",X"03",X"07",X"0F",X"2D",X"2D",X"78",X"2D",X"00",X"00",X"00",X"04",X"06",X"06",X"07",X"07",
		X"00",X"00",X"00",X"08",X"08",X"0C",X"0C",X"0C",X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"2D",X"78",X"2D",X"3C",X"0F",X"07",X"03",X"00",X"07",X"07",X"06",X"06",X"04",X"00",X"00",X"00",
		X"0C",X"0C",X"0C",X"08",X"08",X"00",X"00",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"0F",X"0E",X"00",
		X"22",X"C4",X"48",X"BF",X"48",X"E4",X"B2",X"11",X"99",X"D5",X"72",X"30",X"63",X"F6",X"BB",X"11",
		X"EE",X"AA",X"FF",X"AA",X"AA",X"FF",X"AA",X"AA",X"22",X"22",X"77",X"22",X"22",X"77",X"22",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"77",X"77",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"77",X"00",X"77",X"77",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",
		X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",
		X"00",X"77",X"77",X"77",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"77",X"77",X"00",X"77",
		X"00",X"00",X"00",X"00",X"33",X"74",X"F8",X"F8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"74",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"DD",X"DD",X"DD",X"DD",
		X"00",X"DD",X"DD",X"DD",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"77",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"66",X"66",X"66",X"EE",X"6E",X"08",X"08",X"00",X"00",X"00",X"04",X"06",X"06",X"07",X"07",
		X"00",X"03",X"07",X"0F",X"0D",X"2D",X"78",X"2D",X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"08",X"08",X"4C",X"4C",X"44",X"EE",X"EE",X"00",X"07",X"07",X"06",X"06",X"04",X"00",X"00",X"00",
		X"2D",X"78",X"2D",X"3C",X"0F",X"07",X"03",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"3F",X"3F",X"00",
		X"00",X"EE",X"EE",X"4C",X"4C",X"4C",X"08",X"08",X"00",X"00",X"00",X"04",X"06",X"06",X"07",X"07",
		X"00",X"03",X"07",X"0F",X"2D",X"2D",X"78",X"2D",X"00",X"3F",X"3F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"08",X"08",X"6E",X"EE",X"66",X"66",X"66",X"00",X"07",X"07",X"06",X"06",X"04",X"00",X"00",X"00",
		X"2D",X"78",X"2D",X"3C",X"0F",X"07",X"03",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"0F",X"0E",X"00",
		X"00",X"22",X"22",X"6E",X"6E",X"08",X"08",X"00",X"EE",X"33",X"EE",X"00",X"00",X"11",X"11",X"11",
		X"00",X"FF",X"11",X"77",X"EF",X"CF",X"DF",X"FF",X"00",X"CC",X"CF",X"9E",X"BC",X"AD",X"AD",X"AD",
		X"00",X"08",X"08",X"6E",X"6E",X"22",X"22",X"00",X"11",X"11",X"11",X"00",X"00",X"EE",X"33",X"EE",
		X"FF",X"DF",X"CF",X"EF",X"77",X"11",X"FF",X"00",X"AD",X"AD",X"AD",X"BC",X"9E",X"CF",X"CC",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"88",X"08",X"08",X"00",X"00",X"11",X"33",X"33",X"77",X"77",X"77",
		X"00",X"77",X"FF",X"FF",X"FF",X"BF",X"BF",X"FF",X"00",X"CC",X"EE",X"FF",X"FF",X"FF",X"8F",X"BC",
		X"08",X"08",X"88",X"EE",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"33",X"33",X"11",X"00",X"00",
		X"FF",X"BF",X"BF",X"FF",X"FF",X"FF",X"77",X"00",X"BC",X"8F",X"FF",X"FF",X"FF",X"EE",X"CC",X"00",
		X"00",X"20",X"A0",X"A0",X"A0",X"E0",X"E0",X"A4",X"00",X"00",X"22",X"11",X"00",X"00",X"66",X"00",
		X"00",X"44",X"44",X"00",X"66",X"FF",X"FF",X"FF",X"00",X"00",X"30",X"70",X"F1",X"F3",X"F2",X"F0",
		X"A4",X"E0",X"E0",X"A0",X"A0",X"A0",X"20",X"00",X"00",X"22",X"44",X"00",X"11",X"00",X"00",X"00",
		X"66",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"F0",X"F2",X"73",X"71",X"70",X"30",X"00",X"00",
		X"00",X"02",X"0A",X"0A",X"0A",X"0E",X"0E",X"4A",X"00",X"00",X"22",X"11",X"00",X"00",X"66",X"00",
		X"00",X"44",X"44",X"00",X"66",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"07",X"1E",X"3C",X"2D",X"0F",
		X"4A",X"0E",X"0E",X"0A",X"0A",X"0A",X"02",X"00",X"00",X"22",X"44",X"00",X"11",X"00",X"00",X"00",
		X"66",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"0F",X"2D",X"34",X"16",X"07",X"03",X"00",X"00",
		X"00",X"02",X"0A",X"0A",X"0A",X"0E",X"0E",X"4E",X"00",X"00",X"22",X"11",X"00",X"00",X"66",X"00",
		X"00",X"44",X"44",X"00",X"66",X"FF",X"FF",X"FF",X"00",X"00",X"03",X"07",X"0E",X"0C",X"0D",X"0F",
		X"4E",X"0E",X"0E",X"0A",X"0A",X"0A",X"02",X"00",X"00",X"22",X"44",X"00",X"11",X"00",X"00",X"00",
		X"66",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"0F",X"0D",X"04",X"06",X"07",X"03",X"00",X"00",
		X"66",X"22",X"0E",X"4A",X"C2",X"86",X"84",X"84",X"00",X"00",X"22",X"11",X"00",X"00",X"66",X"00",
		X"00",X"44",X"44",X"00",X"66",X"FF",X"FF",X"FF",X"00",X"00",X"33",X"67",X"AF",X"AF",X"AF",X"EF",
		X"84",X"84",X"86",X"C2",X"4A",X"0E",X"22",X"66",X"00",X"22",X"44",X"00",X"11",X"00",X"00",X"00",
		X"66",X"00",X"00",X"88",X"00",X"00",X"00",X"00",X"EF",X"AF",X"AF",X"AF",X"67",X"33",X"00",X"00",
		X"00",X"00",X"00",X"08",X"3F",X"3F",X"08",X"08",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"74",
		X"00",X"03",X"8F",X"8F",X"AD",X"AD",X"F8",X"AD",X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"08",X"08",X"3F",X"3F",X"08",X"00",X"00",X"00",X"74",X"77",X"33",X"33",X"33",X"11",X"00",X"00",
		X"AD",X"F8",X"AD",X"BC",X"8F",X"8F",X"03",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"0F",X"0E",X"00",
		X"00",X"33",X"33",X"3B",X"3F",X"3F",X"08",X"08",X"00",X"00",X"11",X"33",X"33",X"33",X"77",X"74",
		X"00",X"03",X"8F",X"8F",X"AD",X"AD",X"F8",X"AD",X"00",X"0E",X"0F",X"0F",X"E1",X"A5",X"F0",X"A5",
		X"08",X"08",X"3F",X"3F",X"3B",X"33",X"33",X"00",X"74",X"77",X"33",X"33",X"33",X"11",X"00",X"00",
		X"AD",X"F8",X"AD",X"BC",X"8F",X"8F",X"03",X"00",X"A5",X"F0",X"A5",X"A5",X"0F",X"0F",X"0E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"33",X"77",X"FF",X"FF",X"EF",X"EF",
		X"3F",X"3F",X"BF",X"FF",X"FF",X"FF",X"FF",X"FF",X"10",X"10",X"10",X"30",X"30",X"21",X"30",X"30",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"1E",X"3C",X"F0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"77",X"77",X"11",X"11",X"DD",X"DD",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FC",X"FC",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"F3",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"BF",X"3F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"FF",X"FF",X"EF",X"EF",X"FF",X"FF",X"77",
		X"FF",X"FF",X"77",X"FF",X"FF",X"00",X"00",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"EE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"EE",X"33",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",
		X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"DD",X"DD",X"11",X"11",X"77",
		X"CC",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"77",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"1F",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",
		X"00",X"00",X"00",X"F0",X"F0",X"F0",X"F0",X"F0",X"00",X"00",X"33",X"77",X"FF",X"FF",X"8F",X"8F",
		X"1F",X"1F",X"1F",X"9F",X"FF",X"FF",X"FF",X"9F",X"10",X"10",X"10",X"30",X"30",X"21",X"30",X"30",
		X"F0",X"F0",X"F0",X"F0",X"3C",X"1E",X"3C",X"F0",X"CF",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"FF",X"FF",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"00",X"CC",X"EE",X"F3",X"F3",X"F3",X"F3",X"F3",X"00",X"00",X"00",X"00",X"00",X"88",X"CC",X"EE",
		X"66",X"EE",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"FF",X"FF",X"FF",X"DD",X"CC",X"CC",X"CC",X"DD",
		X"1F",X"1F",X"1F",X"1F",X"1F",X"FF",X"FF",X"FF",X"10",X"10",X"10",X"10",X"10",X"10",X"00",X"00",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"FF",X"EF",X"CF",X"8F",X"8F",X"FF",X"FF",X"77",
		X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"66",X"66",X"00",X"00",X"00",X"00",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"F3",X"FF",X"FF",X"FF",X"EE",X"CC",X"88",X"00",X"00",
		X"CC",X"EE",X"EE",X"EE",X"EE",X"EE",X"EE",X"CC",X"FF",X"FF",X"EE",X"FF",X"FF",X"00",X"00",X"00",
		X"EE",X"DD",X"11",X"FF",X"FF",X"11",X"11",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"33",
		X"00",X"00",X"11",X"77",X"FF",X"FF",X"FF",X"FF",X"00",X"77",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"CF",X"CF",X"CF",X"CF",X"CF",X"33",X"33",X"33",X"77",X"77",X"77",X"77",X"77",
		X"FF",X"0F",X"9E",X"DE",X"FF",X"FF",X"FF",X"FF",X"FF",X"1F",X"F1",X"F1",X"1F",X"9F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"CC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"CC",X"EE",X"EE",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"0F",X"0F",X"0F",X"8F",X"8F",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",
		X"CF",X"CF",X"CF",X"CF",X"CF",X"FF",X"FF",X"FF",X"77",X"77",X"77",X"77",X"77",X"33",X"33",X"33",
		X"FF",X"FF",X"FF",X"FF",X"DE",X"9E",X"0F",X"FF",X"FF",X"FF",X"9F",X"1F",X"F1",X"F1",X"1F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"33",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"77",X"11",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"7F",X"7F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",
		X"8F",X"8F",X"0F",X"0F",X"0F",X"FF",X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"CC",X"00",
		X"FF",X"FF",X"EE",X"EE",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"CF",X"CF",X"CF",X"CF",X"CF",X"FC",X"CF",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"33",
		X"00",X"00",X"11",X"77",X"FF",X"CF",X"CF",X"9E",X"00",X"77",X"FF",X"FF",X"FF",X"0F",X"0F",X"F0",
		X"CF",X"CF",X"CF",X"CF",X"FC",X"CF",X"CF",X"CF",X"33",X"33",X"33",X"33",X"77",X"77",X"77",X"77",
		X"9E",X"9E",X"9E",X"9E",X"CF",X"CF",X"FF",X"FF",X"F0",X"F0",X"F0",X"F0",X"0F",X"0F",X"FF",X"FF",
		X"00",X"00",X"00",X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"2D",X"2D",X"2D",X"2D",X"2D",X"F0",X"2D",
		X"00",X"1F",X"1F",X"1F",X"1F",X"1F",X"F1",X"1F",X"00",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",
		X"EE",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"2D",X"2D",X"2D",X"F0",X"2D",X"2D",X"2D",
		X"1F",X"1F",X"1F",X"1F",X"F1",X"1F",X"1F",X"1F",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"88",
		X"CF",X"CF",X"CF",X"FC",X"CF",X"CF",X"CF",X"CF",X"77",X"77",X"77",X"77",X"33",X"33",X"33",X"33",
		X"FF",X"FF",X"CF",X"CF",X"9E",X"9E",X"9E",X"9E",X"FF",X"FF",X"0F",X"0F",X"F0",X"F0",X"F0",X"F0",
		X"CF",X"FC",X"CF",X"CF",X"CF",X"CF",X"CF",X"00",X"33",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"9E",X"CF",X"CF",X"FF",X"77",X"11",X"00",X"00",X"F0",X"0F",X"0F",X"FF",X"FF",X"FF",X"77",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"2D",X"2D",X"2D",X"F0",X"2D",X"2D",X"2D",X"2D",
		X"1F",X"1F",X"1F",X"F1",X"1F",X"1F",X"1F",X"1F",X"88",X"88",X"88",X"88",X"88",X"88",X"FF",X"FF",
		X"EE",X"EE",X"EE",X"EE",X"EE",X"00",X"00",X"00",X"2D",X"F0",X"2D",X"2D",X"2D",X"2D",X"2D",X"00",
		X"1F",X"F1",X"1F",X"1F",X"1F",X"1F",X"1F",X"00",X"FF",X"FF",X"88",X"88",X"88",X"88",X"88",X"00",
		X"00",X"AA",X"AA",X"EE",X"EE",X"88",X"88",X"88",X"00",X"00",X"11",X"33",X"23",X"67",X"77",X"77",
		X"00",X"67",X"EF",X"3E",X"E3",X"E3",X"3E",X"EF",X"00",X"4B",X"4B",X"F0",X"4B",X"4B",X"F0",X"4B",
		X"88",X"88",X"88",X"EE",X"EE",X"AA",X"AA",X"00",X"77",X"77",X"67",X"23",X"33",X"11",X"00",X"00",
		X"EF",X"3E",X"E3",X"E3",X"3E",X"EF",X"67",X"00",X"4B",X"F0",X"4B",X"4B",X"F0",X"4B",X"4B",X"00",
		X"00",X"00",X"00",X"00",X"EE",X"08",X"08",X"08",X"00",X"00",X"11",X"33",X"23",X"77",X"77",X"77",
		X"00",X"77",X"FF",X"FF",X"3F",X"E3",X"AF",X"EF",X"00",X"CC",X"EE",X"FF",X"FF",X"0F",X"0F",X"6F",
		X"08",X"08",X"08",X"EE",X"00",X"00",X"00",X"00",X"77",X"77",X"77",X"23",X"33",X"11",X"00",X"00",
		X"EF",X"AF",X"E3",X"3F",X"FF",X"FF",X"77",X"00",X"6F",X"0F",X"0F",X"FF",X"FF",X"EE",X"CC",X"00",
		X"00",X"66",X"66",X"66",X"E6",X"E6",X"08",X"08",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"70",X"F0",X"F0",X"F0",X"F7",X"F7",X"F2",X"00",X"C0",X"E0",X"F0",X"F0",X"F0",X"87",X"B4",
		X"08",X"08",X"C0",X"C0",X"40",X"EE",X"EE",X"00",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",
		X"F2",X"F7",X"F7",X"F0",X"F0",X"F0",X"70",X"00",X"B4",X"87",X"F0",X"F0",X"F0",X"F3",X"F3",X"00",
		X"00",X"EE",X"EE",X"40",X"48",X"48",X"08",X"08",X"00",X"00",X"10",X"30",X"30",X"70",X"70",X"70",
		X"00",X"70",X"F0",X"F0",X"F0",X"F7",X"F7",X"F2",X"00",X"F3",X"F3",X"F0",X"87",X"B4",X"B4",X"B4",
		X"08",X"08",X"6E",X"6E",X"66",X"66",X"00",X"00",X"70",X"70",X"70",X"30",X"30",X"10",X"00",X"00",
		X"F2",X"F7",X"F7",X"F0",X"F0",X"F0",X"70",X"00",X"B4",X"B4",X"B4",X"87",X"F0",X"E0",X"C0",X"00",
		X"00",X"66",X"66",X"66",X"6E",X"6E",X"80",X"80",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",
		X"00",X"07",X"0F",X"0F",X"FF",X"F8",X"F8",X"FD",X"00",X"0C",X"0E",X"0F",X"8F",X"8F",X"F8",X"CB",
		X"80",X"80",X"4C",X"4C",X"04",X"EE",X"EE",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",
		X"FD",X"F8",X"F8",X"FF",X"0F",X"0F",X"07",X"00",X"CB",X"F8",X"8F",X"8F",X"0F",X"3F",X"3F",X"00",
		X"00",X"EE",X"EE",X"04",X"0C",X"0C",X"80",X"80",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",
		X"00",X"07",X"0F",X"0F",X"FF",X"F8",X"F8",X"FD",X"00",X"3F",X"3F",X"0F",X"8F",X"8F",X"F8",X"CB",
		X"80",X"80",X"6E",X"6E",X"66",X"66",X"66",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",
		X"FD",X"F8",X"F8",X"FF",X"0F",X"0F",X"07",X"00",X"CB",X"F8",X"8F",X"8F",X"0F",X"0E",X"0C",X"00",
		X"00",X"66",X"66",X"66",X"E6",X"E6",X"80",X"80",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",
		X"00",X"07",X"0F",X"0F",X"0F",X"08",X"08",X"0D",X"00",X"0C",X"0E",X"3C",X"78",X"78",X"78",X"7B",
		X"80",X"80",X"84",X"84",X"04",X"EE",X"EE",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",
		X"0D",X"08",X"08",X"0F",X"0F",X"0F",X"07",X"00",X"7B",X"78",X"78",X"78",X"3C",X"3F",X"3F",X"00",
		X"00",X"EE",X"EE",X"04",X"84",X"84",X"80",X"80",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"07",
		X"00",X"07",X"0F",X"0F",X"0F",X"08",X"08",X"0D",X"00",X"3F",X"3F",X"3C",X"78",X"78",X"78",X"7B",
		X"80",X"80",X"E6",X"E6",X"66",X"66",X"66",X"00",X"07",X"07",X"07",X"03",X"03",X"01",X"00",X"00",
		X"0D",X"08",X"08",X"0F",X"0F",X"0F",X"07",X"00",X"7B",X"78",X"78",X"78",X"3C",X"0E",X"0C",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"08",X"08",X"06",X"02",X"0C",X"00",X"02",X"02",X"0A",X"06",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"00",X"0F",X"04",X"02",X"01",X"02",X"0C",X"00",X"08",X"0E",X"08",X"08",X"08",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"00",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"07",X"00",X"06",X"09",X"09",X"09",X"06",X"02",X"0C",X"00",X"0C",X"02",X"02",X"02",X"0C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"08",X"08",X"07",X"00",X"07",X"08",X"08",X"0C",X"02",X"02",X"0C",X"00",X"0C",X"02",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0C",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"88",X"EE",X"88",X"88",X"88",X"00",X"30",X"70",X"70",X"70",X"F0",X"96",X"96",
		X"00",X"77",X"FF",X"FF",X"9F",X"9F",X"FF",X"FF",X"00",X"EE",X"FF",X"FF",X"FF",X"FF",X"F9",X"F9",
		X"88",X"EE",X"88",X"00",X"00",X"00",X"00",X"00",X"F0",X"70",X"70",X"70",X"30",X"77",X"77",X"77",
		X"9F",X"9F",X"FF",X"FF",X"77",X"11",X"FF",X"00",X"FF",X"FF",X"FF",X"FF",X"EE",X"00",X"00",X"00",
		X"00",X"22",X"AA",X"EE",X"EE",X"88",X"88",X"88",X"00",X"30",X"70",X"70",X"70",X"F0",X"96",X"96",
		X"00",X"77",X"FF",X"8F",X"CF",X"EF",X"FF",X"FF",X"00",X"EE",X"FF",X"F8",X"F8",X"F8",X"F8",X"F8",
		X"88",X"EE",X"EE",X"AA",X"22",X"CC",X"CC",X"CC",X"F0",X"70",X"70",X"70",X"30",X"00",X"00",X"00",
		X"EF",X"CF",X"8F",X"FF",X"77",X"11",X"00",X"00",X"F8",X"F8",X"F8",X"FF",X"EE",X"99",X"FF",X"11",
		X"00",X"22",X"22",X"22",X"66",X"CC",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"21",
		X"00",X"00",X"D1",X"F3",X"F3",X"E3",X"E3",X"7B",X"00",X"EE",X"FF",X"FD",X"FD",X"FD",X"FD",X"FD",
		X"00",X"00",X"CC",X"66",X"22",X"22",X"22",X"00",X"21",X"30",X"10",X"10",X"10",X"00",X"00",X"00",
		X"7B",X"E3",X"E3",X"F3",X"F3",X"D1",X"00",X"00",X"FD",X"FD",X"FD",X"FD",X"FD",X"FF",X"EE",X"00",
		X"00",X"66",X"AA",X"EE",X"E6",X"E6",X"E6",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"30",X"70",X"70",X"70",X"F0",X"96",X"00",X"33",X"77",X"FF",X"DF",X"9F",X"BF",X"FF",
		X"E6",X"E6",X"E6",X"E6",X"EE",X"AA",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"96",X"F0",X"70",X"70",X"70",X"30",X"00",X"00",X"FF",X"BF",X"9F",X"DF",X"FF",X"77",X"33",X"00",
		X"00",X"66",X"22",X"AA",X"EE",X"E6",X"E6",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"21",X"00",X"00",X"C0",X"D1",X"F3",X"F3",X"F3",X"7B",
		X"E6",X"E6",X"E6",X"EE",X"AA",X"22",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"30",X"10",X"10",X"10",X"00",X"00",X"00",X"7B",X"F3",X"F3",X"F3",X"D1",X"C0",X"00",X"00",
		X"00",X"66",X"22",X"22",X"EE",X"EA",X"EA",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"70",X"70",X"70",X"F0",X"96",
		X"EA",X"EA",X"EA",X"EE",X"22",X"22",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"F0",X"70",X"70",X"70",X"30",X"00",X"00",
		X"00",X"00",X"60",X"E0",X"E0",X"E0",X"E0",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",
		X"2C",X"E0",X"E0",X"E0",X"E0",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"44",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"70",X"70",X"70",X"F0",X"96",
		X"00",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"96",X"F0",X"70",X"70",X"70",X"30",X"00",X"00",
		X"00",X"00",X"00",X"22",X"22",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"10",X"10",X"30",X"21",X"00",X"00",X"C0",X"C0",X"C0",X"F3",X"C0",X"48",
		X"00",X"00",X"EE",X"22",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"21",X"30",X"10",X"10",X"10",X"00",X"00",X"00",X"48",X"C0",X"F3",X"C0",X"C0",X"C0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"44",X"11",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"11",X"00",X"00",X"00",X"11",X"99",X"44",X"00",X"00",
		X"00",X"22",X"11",X"88",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"22",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"88",X"22",X"22",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
