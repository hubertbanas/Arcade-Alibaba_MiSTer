library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ROM_PGM_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ROM_PGM_1 is
	type rom is array(0 to  10239) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"01",X"03",X"04",X"02",X"01",X"03",X"02",X"04",X"02",X"03",X"04",X"01",X"01",X"02",X"04",X"03",
		X"02",X"03",X"01",X"04",X"03",X"02",X"04",X"01",X"01",X"01",X"03",X"04",X"02",X"01",X"04",X"03",
		X"03",X"02",X"01",X"04",X"04",X"02",X"03",X"01",X"02",X"01",X"03",X"04",X"03",X"01",X"04",X"02",
		X"04",X"02",X"01",X"03",X"03",X"01",X"02",X"04",X"04",X"01",X"03",X"02",X"04",X"01",X"02",X"03",
		X"00",X"04",X"08",X"0C",X"10",X"14",X"18",X"1C",X"20",X"24",X"28",X"2C",X"30",X"34",X"38",X"3C",
		X"F5",X"E5",X"D5",X"3A",X"C0",X"50",X"E6",X"0F",X"5F",X"16",X"00",X"21",X"40",X"80",X"19",X"5E",
		X"21",X"00",X"80",X"19",X"11",X"E0",X"4D",X"01",X"04",X"00",X"ED",X"B0",X"D1",X"E1",X"F1",X"C9",
		X"F5",X"AF",X"32",X"80",X"50",X"00",X"00",X"00",X"F1",X"C9",X"CD",X"0F",X"20",X"FE",X"FC",X"28",
		X"02",X"FE",X"FD",X"CA",X"40",X"19",X"FE",X"70",X"C3",X"F0",X"88",X"7D",X"21",X"E0",X"4D",X"FE",
		X"EB",X"28",X"14",X"FE",X"90",X"20",X"03",X"23",X"18",X"0D",X"FE",X"F4",X"20",X"04",X"23",X"23",
		X"18",X"05",X"FE",X"70",X"23",X"23",X"23",X"7E",X"32",X"E4",X"4D",X"3E",X"72",X"CD",X"9E",X"3E",
		X"3E",X"11",X"CD",X"AB",X"3E",X"C3",X"75",X"8E",X"FF",X"FF",X"FF",X"3A",X"E6",X"4D",X"A7",X"C0",
		X"3E",X"01",X"32",X"E6",X"4D",X"CD",X"3D",X"81",X"CD",X"2D",X"83",X"C9",X"3E",X"01",X"06",X"03",
		X"11",X"20",X"00",X"C5",X"D5",X"E5",X"CF",X"E1",X"D1",X"C1",X"C9",X"21",X"CD",X"45",X"CD",X"CC",
		X"80",X"19",X"CD",X"CC",X"80",X"19",X"CD",X"CC",X"80",X"19",X"CD",X"CC",X"80",X"C9",X"01",X"FD",
		X"80",X"21",X"D0",X"41",X"CD",X"72",X"81",X"3E",X"DA",X"32",X"30",X"42",X"C9",X"DA",X"DA",X"DA",
		X"CD",X"69",X"8B",X"CD",X"77",X"8D",X"CD",X"DB",X"80",X"CD",X"EE",X"80",X"C9",X"00",X"00",X"00",
		X"3A",X"1C",X"4E",X"C6",X"99",X"27",X"CD",X"A8",X"85",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"C6",
		X"30",X"32",X"F2",X"41",X"3A",X"1C",X"4E",X"E6",X"0F",X"C6",X"30",X"32",X"D2",X"41",X"3E",X"0F",
		X"32",X"F2",X"45",X"32",X"D2",X"45",X"CD",X"B2",X"82",X"C9",X"F0",X"72",X"F1",X"3E",X"11",X"CD",
		X"99",X"0F",X"01",X"3A",X"81",X"21",X"84",X"40",X"CD",X"72",X"81",X"21",X"64",X"41",X"CD",X"72",
		X"81",X"21",X"44",X"42",X"CD",X"72",X"81",X"21",X"24",X"43",X"CD",X"72",X"81",X"C9",X"3E",X"17",
		X"CD",X"99",X"0F",X"01",X"ED",X"0F",X"CD",X"45",X"81",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C5",X"00",X"11",X"20",X"00",X"0A",X"77",X"19",X"03",X"0A",X"77",X"19",X"03",X"0A",
		X"77",X"C1",X"C9",X"3A",X"FA",X"4D",X"A7",X"C0",X"3A",X"E6",X"4D",X"A7",X"C0",X"3E",X"01",X"32",
		X"E6",X"4D",X"CD",X"3D",X"81",X"CD",X"2D",X"83",X"21",X"9C",X"4E",X"36",X"10",X"C9",X"21",X"BC",
		X"4E",X"36",X"02",X"21",X"04",X"4E",X"C9",X"21",X"90",X"4C",X"3A",X"8A",X"4C",X"4F",X"06",X"10",
		X"7E",X"A7",X"28",X"2F",X"E6",X"C0",X"07",X"07",X"B9",X"30",X"28",X"35",X"7E",X"E6",X"3F",X"20",
		X"22",X"77",X"C5",X"E5",X"2C",X"7E",X"2C",X"46",X"21",X"E1",X"81",X"E5",X"E7",X"94",X"08",X"A3",
		X"06",X"8E",X"05",X"42",X"12",X"00",X"10",X"0B",X"10",X"63",X"02",X"2B",X"21",X"F0",X"21",X"B9",
		X"22",X"E1",X"C1",X"2C",X"2C",X"2C",X"10",X"C8",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3A",X"ED",X"4D",X"A7",X"20",X"09",X"3E",X"01",X"32",X"ED",X"4D",X"CD",X"E9",
		X"0F",X"C9",X"3A",X"EF",X"4D",X"A7",X"20",X"04",X"CD",X"79",X"3F",X"C9",X"C3",X"61",X"84",X"00",
		X"21",X"00",X"40",X"CF",X"06",X"3F",X"21",X"C0",X"43",X"CF",X"3A",X"EE",X"4D",X"A7",X"C0",X"3E",
		X"01",X"32",X"E8",X"4D",X"CD",X"82",X"3C",X"C9",X"3A",X"E8",X"4D",X"A7",X"C0",X"3A",X"09",X"4E",
		X"C3",X"47",X"03",X"CD",X"3E",X"75",X"21",X"37",X"43",X"11",X"20",X"00",X"77",X"3D",X"19",X"77",
		X"3E",X"05",X"32",X"37",X"47",X"32",X"57",X"47",X"CD",X"8A",X"05",X"C9",X"1F",X"C9",X"AF",X"32",
		X"B1",X"4D",X"C9",X"F1",X"02",X"F2",X"03",X"F3",X"0F",X"70",X"F4",X"02",X"8D",X"F4",X"02",X"88",
		X"F4",X"02",X"8A",X"70",X"F4",X"01",X"6C",X"F4",X"02",X"8A",X"F4",X"01",X"6A",X"F4",X"02",X"88",
		X"70",X"F4",X"02",X"8D",X"F4",X"02",X"88",X"F4",X"02",X"8A",X"70",X"F4",X"01",X"6C",X"F4",X"02",
		X"8A",X"F4",X"01",X"6A",X"F4",X"02",X"88",X"70",X"F0",X"6A",X"82",X"FF",X"21",X"BC",X"4E",X"CB",
		X"AE",X"3E",X"01",X"32",X"F5",X"90",X"C9",X"3E",X"01",X"32",X"F4",X"90",X"CD",X"9C",X"82",X"CB",
		X"F6",X"C9",X"3A",X"EA",X"90",X"A7",X"C0",X"CD",X"00",X"8F",X"C9",X"3E",X"01",X"32",X"80",X"50",
		X"C9",X"3E",X"00",X"32",X"80",X"50",X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"28",X"10",X"AF",X"32",
		X"80",X"50",X"CD",X"51",X"8C",X"CD",X"00",X"81",X"3E",X"02",X"32",X"80",X"50",X"C9",X"3A",X"1C",
		X"4E",X"A7",X"20",X"10",X"CD",X"C0",X"8C",X"3A",X"FB",X"4D",X"21",X"16",X"4E",X"86",X"77",X"3E",
		X"40",X"32",X"1C",X"4E",X"AF",X"21",X"E0",X"4D",X"06",X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",
		X"CF",X"CD",X"00",X"81",X"CD",X"35",X"A4",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",
		X"00",X"00",X"22",X"FC",X"4D",X"22",X"FE",X"4D",X"C9",X"CD",X"7C",X"0E",X"3E",X"20",X"32",X"04",
		X"4E",X"C9",X"CD",X"6C",X"0E",X"CD",X"B0",X"0E",X"CD",X"C1",X"2C",X"C9",X"FF",X"06",X"16",X"CD",
		X"5E",X"2C",X"C9",X"FF",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"08",X"DD",X"21",X"E9",X"4D",X"C9",
		X"DD",X"21",X"39",X"4D",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"06",X"3A",X"AF",X"4D",X"C3",
		X"4C",X"3D",X"3A",X"AC",X"4D",X"A7",X"28",X"06",X"3A",X"AF",X"4D",X"C3",X"4C",X"3D",X"3A",X"F9",
		X"4D",X"A7",X"C2",X"83",X"83",X"3A",X"16",X"4E",X"A7",X"CA",X"4C",X"83",X"2A",X"31",X"4D",X"11",
		X"22",X"23",X"A7",X"ED",X"52",X"C2",X"4C",X"83",X"3E",X"08",X"32",X"F9",X"4D",X"C3",X"4C",X"83",
		X"00",X"00",X"00",X"2A",X"31",X"4D",X"11",X"3A",X"2D",X"A7",X"ED",X"52",X"C2",X"4C",X"83",X"AF",
		X"32",X"F9",X"4D",X"C3",X"45",X"83",X"00",X"00",X"00",X"3A",X"E4",X"4D",X"FE",X"01",X"C2",X"02",
		X"3E",X"3E",X"01",X"32",X"A7",X"4D",X"C3",X"63",X"17",X"2A",X"39",X"4D",X"7D",X"06",X"23",X"90",
		X"3A",X"39",X"4D",X"D8",X"06",X"25",X"90",X"D8",X"CD",X"D6",X"A0",X"C9",X"FF",X"FF",X"CD",X"FB",
		X"83",X"21",X"00",X"00",X"28",X"03",X"22",X"FC",X"4D",X"22",X"FE",X"4D",X"C9",X"00",X"00",X"00",
		X"00",X"E5",X"D5",X"11",X"20",X"00",X"77",X"3C",X"19",X"77",X"3C",X"3C",X"23",X"77",X"3D",X"ED",
		X"52",X"77",X"D1",X"E1",X"C9",X"CD",X"17",X"2D",X"3A",X"00",X"4E",X"FE",X"03",X"D0",X"CD",X"F3",
		X"2C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"E4",X"4D",X"FE",X"01",
		X"C9",X"FD",X"21",X"0A",X"4D",X"CD",X"FB",X"83",X"28",X"09",X"DD",X"21",X"E9",X"4D",X"CD",X"FA",
		X"09",X"18",X"03",X"CD",X"A9",X"31",X"30",X"0E",X"3A",X"B1",X"4D",X"A7",X"C0",X"3E",X"01",X"32",
		X"B1",X"4D",X"CD",X"07",X"1F",X"C9",X"AF",X"32",X"B1",X"4D",X"C9",X"F5",X"E5",X"D5",X"11",X"00",
		X"04",X"3E",X"11",X"19",X"77",X"D1",X"E1",X"F1",X"77",X"C9",X"D5",X"E5",X"06",X"20",X"4F",X"CD",
		X"2B",X"84",X"F5",X"E5",X"11",X"E0",X"83",X"7D",X"E6",X"1F",X"87",X"26",X"00",X"6F",X"19",X"D1",
		X"A7",X"ED",X"52",X"F1",X"EE",X"01",X"CD",X"2B",X"84",X"EB",X"23",X"79",X"10",X"E1",X"E1",X"D1",
		X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"C2",X"2A",X"82",X"3E",X"40",X"06",X"3F",X"C3",X"20",X"82",
		X"2A",X"B0",X"8F",X"22",X"86",X"4D",X"11",X"B2",X"8F",X"01",X"20",X"00",X"1A",X"FE",X"FF",X"C8",
		X"FE",X"FE",X"20",X"0A",X"2A",X"86",X"4D",X"23",X"22",X"86",X"4D",X"13",X"18",X"EE",X"77",X"E5",
		X"C5",X"01",X"00",X"04",X"09",X"3E",X"01",X"77",X"C1",X"E1",X"09",X"13",X"18",X"DE",X"2A",X"24",
		X"4C",X"ED",X"5B",X"26",X"4C",X"ED",X"4B",X"28",X"4C",X"22",X"26",X"4C",X"ED",X"53",X"28",X"4C",
		X"2A",X"2A",X"4C",X"ED",X"43",X"2A",X"4C",X"22",X"24",X"4C",X"2A",X"34",X"4C",X"ED",X"5B",X"36",
		X"4C",X"ED",X"4B",X"38",X"4C",X"22",X"36",X"4C",X"ED",X"53",X"38",X"4C",X"2A",X"3A",X"4C",X"ED",
		X"43",X"3A",X"4C",X"22",X"34",X"4C",X"C9",X"21",X"83",X"E3",X"22",X"02",X"4D",X"21",X"83",X"D1",
		X"22",X"04",X"4D",X"21",X"83",X"BF",X"22",X"06",X"4D",X"CD",X"99",X"14",X"C9",X"21",X"97",X"D1",
		X"22",X"00",X"4D",X"CD",X"99",X"14",X"C9",X"3E",X"94",X"21",X"34",X"43",X"77",X"E5",X"23",X"3C",
		X"77",X"23",X"3C",X"77",X"E1",X"11",X"20",X"00",X"19",X"3C",X"77",X"23",X"3C",X"77",X"23",X"3C",
		X"77",X"3E",X"01",X"21",X"34",X"47",X"11",X"20",X"00",X"01",X"00",X"03",X"E5",X"C5",X"CF",X"C1",
		X"E1",X"19",X"CF",X"C9",X"3E",X"01",X"CD",X"74",X"0F",X"C9",X"01",X"5A",X"85",X"CD",X"72",X"81",
		X"C9",X"E5",X"CD",X"2A",X"85",X"E1",X"11",X"00",X"04",X"19",X"CD",X"24",X"85",X"C9",X"21",X"50",
		X"40",X"CD",X"31",X"85",X"C9",X"21",X"53",X"40",X"CD",X"31",X"85",X"C9",X"21",X"55",X"40",X"CD",
		X"31",X"85",X"C9",X"21",X"57",X"40",X"CD",X"31",X"85",X"C9",X"53",X"54",X"50",X"AF",X"32",X"FB",
		X"4D",X"21",X"00",X"00",X"22",X"A4",X"4D",X"21",X"31",X"93",X"22",X"08",X"4D",X"CD",X"99",X"14",
		X"06",X"01",X"CD",X"ED",X"23",X"CD",X"B3",X"85",X"CD",X"8A",X"05",X"C9",X"21",X"FB",X"4D",X"19",
		X"D5",X"E5",X"11",X"A7",X"4D",X"A7",X"ED",X"52",X"E1",X"D1",X"06",X"02",X"28",X"0A",X"06",X"00",
		X"7E",X"A7",X"28",X"07",X"06",X"01",X"AF",X"77",X"CD",X"CD",X"0F",X"CD",X"10",X"81",X"CD",X"5A",
		X"2A",X"CD",X"12",X"86",X"00",X"E6",X"C9",X"C9",X"32",X"1C",X"4E",X"A7",X"C0",X"3E",X"01",X"32",
		X"DF",X"90",X"C9",X"CD",X"70",X"84",X"CD",X"38",X"8E",X"C9",X"FF",X"FF",X"21",X"00",X"00",X"22",
		X"08",X"4D",X"22",X"02",X"4D",X"22",X"04",X"4D",X"22",X"06",X"4D",X"22",X"00",X"4D",X"22",X"F0",
		X"90",X"22",X"F2",X"90",X"22",X"D2",X"4D",X"22",X"E4",X"4D",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",
		X"20",X"04",X"CD",X"56",X"89",X"C9",X"FE",X"02",X"20",X"07",X"CD",X"70",X"8B",X"CD",X"49",X"3D",
		X"C9",X"06",X"04",X"ED",X"5B",X"39",X"4D",X"CD",X"23",X"17",X"CD",X"49",X"3D",X"C9",X"21",X"BC",
		X"4E",X"CB",X"DE",X"CD",X"9C",X"82",X"C9",X"FF",X"FF",X"21",X"BC",X"4E",X"CB",X"D6",X"CD",X"9C",
		X"82",X"C9",X"21",X"BC",X"4E",X"36",X"10",X"CD",X"9C",X"82",X"CD",X"17",X"2D",X"C9",X"FF",X"FF",
		X"CD",X"FB",X"83",X"28",X"07",X"DD",X"21",X"01",X"33",X"C3",X"D6",X"10",X"EF",X"04",X"01",X"AF",
		X"32",X"AC",X"4D",X"32",X"A7",X"4D",X"32",X"F0",X"90",X"C3",X"01",X"11",X"21",X"F0",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"4F",X"1B",X"C3",X"C3",X"10",X"21",X"F1",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"C7",X"1B",X"C3",X"1B",X"11",X"21",X"F2",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"3F",X"1C",X"C3",X"5F",X"11",X"21",X"F3",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"B7",X"1C",X"C3",X"CC",X"11",X"3A",X"E4",X"4D",X"32",
		X"FF",X"90",X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"D0",X"3E",X"02",X"32",X"9C",X"4E",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"21",X"06",X"4C",X"06",X"04",X"1A",X"77",X"23",X"23",X"13",X"05",X"20",
		X"F8",X"C9",X"21",X"07",X"4C",X"3E",X"09",X"06",X"04",X"77",X"23",X"23",X"05",X"20",X"FA",X"C9",
		X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"C9",X"CD",X"3F",X"88",X"11",X"61",X"12",X"A7",
		X"C8",X"11",X"65",X"12",X"C9",X"CD",X"33",X"88",X"11",X"69",X"12",X"A7",X"C8",X"11",X"6D",X"12",
		X"C9",X"CD",X"57",X"88",X"11",X"71",X"12",X"A7",X"C8",X"11",X"75",X"12",X"C9",X"CD",X"4B",X"88",
		X"11",X"79",X"12",X"A7",X"C8",X"11",X"7D",X"12",X"C9",X"CD",X"B0",X"86",X"20",X"22",X"3A",X"30",
		X"4D",X"FE",X"00",X"20",X"04",X"CD",X"C5",X"86",X"C9",X"FE",X"01",X"20",X"04",X"CD",X"B9",X"86",
		X"C9",X"FE",X"02",X"20",X"04",X"CD",X"B9",X"86",X"C9",X"FE",X"03",X"C0",X"CD",X"C5",X"86",X"C9",
		X"3A",X"30",X"4D",X"FE",X"00",X"20",X"04",X"CD",X"DD",X"86",X"C9",X"FE",X"01",X"20",X"04",X"CD",
		X"D1",X"86",X"C9",X"FE",X"02",X"20",X"04",X"CD",X"D1",X"86",X"C9",X"FE",X"03",X"C0",X"CD",X"DD",
		X"86",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"04",X"CD",X"9C",X"16",X"C9",X"CD",X"E9",X"86",
		X"CD",X"94",X"86",X"CD",X"A2",X"86",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"04",X"CD",X"AA",
		X"16",X"C9",X"CD",X"E9",X"86",X"CD",X"94",X"86",X"CD",X"A2",X"86",X"C9",X"21",X"02",X"4C",X"CD",
		X"4E",X"15",X"CD",X"32",X"87",X"CD",X"47",X"87",X"C9",X"21",X"00",X"00",X"22",X"01",X"90",X"22",
		X"03",X"90",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"08",X"FE",X"02",X"28",X"04",X"CD",X"09",
		X"3D",X"C9",X"3A",X"FD",X"4D",X"A7",X"C8",X"CD",X"09",X"3D",X"C9",X"3E",X"40",X"06",X"0C",X"21",
		X"45",X"41",X"CD",X"76",X"0F",X"C9",X"00",X"DD",X"21",X"26",X"4D",X"CD",X"0F",X"20",X"21",X"00",
		X"90",X"FE",X"FC",X"28",X"0D",X"FE",X"FD",X"28",X"09",X"E6",X"C0",X"D6",X"C0",X"20",X"03",X"36",
		X"01",X"C9",X"36",X"00",X"C9",X"0D",X"0C",X"0B",X"0A",X"09",X"6C",X"08",X"07",X"00",X"00",X"06",
		X"2A",X"39",X"4D",X"7D",X"06",X"02",X"80",X"32",X"D2",X"4D",X"7C",X"32",X"D3",X"4D",X"C9",X"1E",
		X"3A",X"3C",X"4D",X"FE",X"00",X"20",X"12",X"FD",X"21",X"35",X"4D",X"CD",X"97",X"87",X"7E",X"A7",
		X"C0",X"FD",X"21",X"37",X"4D",X"CD",X"97",X"87",X"C9",X"FE",X"01",X"20",X"15",X"CD",X"C0",X"87",
		X"FD",X"21",X"D2",X"4D",X"CD",X"97",X"87",X"7E",X"A7",X"C0",X"FD",X"21",X"37",X"4D",X"CD",X"97",
		X"87",X"C9",X"FE",X"02",X"20",X"04",X"CD",X"ED",X"87",X"C9",X"FE",X"03",X"C0",X"CD",X"D7",X"87",
		X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"08",X"CD",X"D0",X"87",X"3A",X"00",X"90",X"A7",X"C0",
		X"FD",X"21",X"39",X"4D",X"C3",X"7A",X"80",X"AF",X"21",X"00",X"90",X"01",X"FF",X"03",X"CF",X"C3",
		X"3E",X"A7",X"00",X"CD",X"69",X"87",X"3E",X"01",X"32",X"01",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",
		X"69",X"87",X"3E",X"01",X"32",X"02",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",X"69",X"87",X"3E",X"01",
		X"32",X"03",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",X"69",X"87",X"3E",X"01",X"32",X"04",X"90",X"3A",
		X"C0",X"4D",X"C9",X"06",X"04",X"2A",X"37",X"4D",X"A7",X"ED",X"52",X"28",X"1C",X"05",X"2A",X"35",
		X"4D",X"A7",X"ED",X"52",X"28",X"13",X"05",X"2A",X"39",X"4D",X"A7",X"ED",X"52",X"28",X"0A",X"05",
		X"2A",X"D2",X"4D",X"A7",X"ED",X"52",X"28",X"01",X"05",X"78",X"C9",X"3A",X"FD",X"4D",X"A7",X"3E",
		X"01",X"28",X"03",X"32",X"FB",X"4D",X"32",X"FF",X"90",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"5B",X"33",X"4D",X"CD",X"63",X"88",X"32",X"06",X"90",X"A7",X"C8",X"3E",X"01",X"32",X"A8",
		X"4D",X"3E",X"02",X"32",X"A4",X"4D",X"C9",X"ED",X"5B",X"31",X"4D",X"CD",X"63",X"88",X"32",X"05",
		X"90",X"A7",X"C8",X"3E",X"01",X"32",X"A7",X"4D",X"32",X"A4",X"4D",X"C9",X"00",X"00",X"00",X"3A",
		X"05",X"90",X"A7",X"28",X"0B",X"AF",X"32",X"A7",X"4D",X"32",X"05",X"90",X"32",X"A4",X"4D",X"C9",
		X"3A",X"06",X"90",X"A7",X"C8",X"AF",X"32",X"A8",X"4D",X"32",X"06",X"90",X"32",X"A4",X"4D",X"C9",
		X"CA",X"8B",X"80",X"FE",X"90",X"CA",X"F5",X"18",X"FE",X"92",X"CA",X"F5",X"18",X"C3",X"EF",X"18",
		X"A7",X"C8",X"47",X"CD",X"B0",X"86",X"20",X"04",X"CD",X"28",X"8F",X"C9",X"CD",X"46",X"8F",X"C9",
		X"31",X"C0",X"4F",X"AF",X"01",X"04",X"00",X"21",X"00",X"90",X"CF",X"0D",X"20",X"FC",X"C3",X"3E",
		X"A7",X"00",X"00",X"00",X"C8",X"78",X"FE",X"02",X"C8",X"FE",X"01",X"C8",X"3E",X"01",X"32",X"A4",
		X"4D",X"CD",X"CF",X"88",X"C9",X"D6",X"C0",X"28",X"0A",X"7E",X"FE",X"90",X"28",X"05",X"FE",X"92",
		X"C2",X"9F",X"29",X"11",X"00",X"04",X"19",X"7E",X"FE",X"16",X"CA",X"0B",X"8B",X"FE",X"17",X"CA",
		X"9F",X"29",X"C3",X"C6",X"29",X"FF",X"3A",X"AC",X"4D",X"A7",X"C0",X"00",X"00",X"CD",X"B7",X"88",
		X"3A",X"05",X"90",X"CD",X"00",X"89",X"A7",X"28",X"09",X"AF",X"32",X"08",X"90",X"06",X"02",X"CD",
		X"9B",X"85",X"CD",X"49",X"3D",X"3A",X"AD",X"4D",X"A7",X"C0",X"00",X"00",X"CD",X"A0",X"88",X"3A",
		X"06",X"90",X"CD",X"00",X"89",X"A7",X"20",X"06",X"CD",X"49",X"3D",X"C9",X"00",X"00",X"3A",X"A4",
		X"4D",X"CD",X"6C",X"17",X"AF",X"32",X"FD",X"4D",X"CD",X"49",X"3D",X"C9",X"00",X"00",X"00",X"00",
		X"21",X"02",X"4C",X"CD",X"4E",X"15",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"07",X"CD",X"32",X"87",
		X"CD",X"47",X"87",X"C9",X"FE",X"02",X"C0",X"CD",X"E0",X"89",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"C9",X"CD",X"C0",X"89",X"ED",X"53",X"02",X"4C",X"ED",
		X"43",X"06",X"4C",X"23",X"CD",X"C0",X"89",X"ED",X"53",X"08",X"4C",X"ED",X"43",X"0C",X"4C",X"C9",
		X"3A",X"E4",X"4D",X"FE",X"02",X"C0",X"CD",X"B0",X"86",X"20",X"10",X"3A",X"C0",X"4D",X"21",X"10",
		X"8A",X"A7",X"20",X"03",X"21",X"18",X"8A",X"CD",X"C8",X"89",X"C9",X"3A",X"C0",X"4D",X"21",X"20",
		X"8A",X"A7",X"20",X"03",X"21",X"28",X"8A",X"CD",X"C8",X"89",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"68",X"01",X"60",X"01",X"64",X"01",X"6C",X"01",X"78",X"01",X"70",X"01",X"74",X"01",X"7C",X"01",
		X"6B",X"01",X"63",X"01",X"67",X"01",X"6F",X"01",X"7B",X"01",X"73",X"01",X"77",X"01",X"7F",X"01",
		X"3E",X"FD",X"21",X"85",X"40",X"06",X"15",X"CF",X"21",X"B9",X"40",X"11",X"20",X"00",X"06",X"18",
		X"77",X"19",X"05",X"20",X"FB",X"21",X"8A",X"42",X"06",X"0A",X"CF",X"00",X"00",X"00",X"00",X"21",
		X"CA",X"41",X"06",X"06",X"77",X"19",X"05",X"20",X"FB",X"21",X"AA",X"41",X"77",X"23",X"77",X"21",
		X"73",X"42",X"77",X"C3",X"50",X"8B",X"AF",X"06",X"5F",X"21",X"8C",X"4E",X"CF",X"C9",X"FF",X"FF",
		X"3E",X"40",X"21",X"A5",X"40",X"06",X"14",X"CF",X"21",X"A9",X"42",X"06",X"0B",X"CF",X"21",X"D8",
		X"40",X"06",X"17",X"77",X"19",X"05",X"20",X"FB",X"21",X"A9",X"41",X"06",X"08",X"77",X"19",X"05",
		X"20",X"FB",X"21",X"89",X"41",X"77",X"23",X"77",X"21",X"6F",X"40",X"77",X"23",X"77",X"C9",X"FF",
		X"84",X"44",X"85",X"44",X"88",X"44",X"8E",X"44",X"91",X"44",X"97",X"44",X"39",X"45",X"99",X"45",
		X"79",X"46",X"D9",X"46",X"99",X"47",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"0B",X"11",X"A0",X"8A",X"1A",X"6F",X"13",X"1A",X"67",X"3E",X"16",X"77",X"13",X"05",X"20",
		X"F4",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"07",X"CD",X"00",X"81",X"CD",X"3D",X"25",X"C9",
		X"FE",X"02",X"C0",X"CD",X"00",X"81",X"CD",X"30",X"8A",X"CD",X"70",X"8A",X"CD",X"C0",X"8A",X"CD",
		X"20",X"8D",X"C9",X"FE",X"90",X"CA",X"23",X"19",X"FE",X"92",X"CA",X"23",X"19",X"E6",X"C0",X"D6",
		X"C0",X"CA",X"23",X"19",X"C3",X"50",X"19",X"FF",X"FF",X"FF",X"FF",X"DD",X"E5",X"FD",X"E5",X"00",
		X"00",X"00",X"00",X"FD",X"21",X"0C",X"4D",X"CD",X"0F",X"20",X"19",X"7E",X"FD",X"E1",X"DD",X"E1",
		X"FE",X"16",X"CA",X"9F",X"29",X"C3",X"C6",X"29",X"3A",X"E4",X"4D",X"21",X"00",X"00",X"FE",X"02",
		X"28",X"07",X"FE",X"01",X"C0",X"22",X"FE",X"4D",X"C9",X"22",X"FE",X"4D",X"AF",X"32",X"FC",X"4D",
		X"C9",X"BC",X"02",X"5C",X"40",X"53",X"45",X"47",X"41",X"40",X"31",X"39",X"38",X"32",X"2F",X"81",
		X"21",X"D2",X"D2",X"22",X"4F",X"40",X"21",X"FC",X"FC",X"22",X"4F",X"43",X"22",X"6F",X"43",X"22",
		X"8F",X"43",X"21",X"D3",X"D3",X"22",X"AF",X"43",X"C9",X"CD",X"A3",X"8E",X"CD",X"7F",X"0F",X"C9",
		X"06",X"05",X"ED",X"5B",X"39",X"4D",X"3A",X"AF",X"4D",X"A7",X"20",X"09",X"2A",X"37",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AE",X"4D",X"A7",X"20",X"09",X"2A",X"35",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AD",X"4D",X"A7",X"20",X"09",X"2A",X"33",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AC",X"4D",X"A7",X"20",X"09",X"2A",X"31",X"4D",X"A7",
		X"ED",X"52",X"C3",X"6C",X"8F",X"05",X"CD",X"CD",X"8D",X"00",X"32",X"A5",X"4D",X"A7",X"C8",X"C3",
		X"80",X"8E",X"CD",X"83",X"8F",X"AF",X"32",X"A5",X"4D",X"3A",X"FD",X"4D",X"A7",X"06",X"00",X"28",
		X"09",X"AF",X"32",X"FD",X"4D",X"CD",X"CD",X"0F",X"06",X"01",X"CD",X"10",X"8F",X"C9",X"21",X"02",
		X"4C",X"11",X"F0",X"90",X"06",X"04",X"1A",X"A7",X"28",X"06",X"FE",X"F0",X"20",X"02",X"36",X"FC",
		X"23",X"23",X"13",X"05",X"20",X"F0",X"C9",X"00",X"DD",X"40",X"07",X"C1",X"40",X"40",X"FF",X"FF",
		X"2A",X"17",X"4E",X"3E",X"40",X"CD",X"F4",X"3C",X"11",X"60",X"00",X"19",X"22",X"17",X"4E",X"C9",
		X"2A",X"17",X"4E",X"11",X"60",X"00",X"ED",X"52",X"22",X"17",X"4E",X"3E",X"90",X"CD",X"DE",X"3C",
		X"3E",X"01",X"CD",X"F4",X"3C",X"C9",X"2A",X"1A",X"4E",X"CD",X"1B",X"8C",X"11",X"60",X"00",X"19",
		X"22",X"1A",X"4E",X"C9",X"2A",X"1A",X"4E",X"11",X"60",X"00",X"ED",X"52",X"3E",X"40",X"CD",X"F4",
		X"3C",X"22",X"1A",X"4E",X"C9",X"21",X"FB",X"4D",X"35",X"21",X"16",X"4E",X"34",X"CD",X"10",X"8C",
		X"C9",X"01",X"0B",X"00",X"CD",X"FA",X"8D",X"11",X"16",X"4E",X"ED",X"B0",X"C9",X"00",X"00",X"00",
		X"00",X"7E",X"A7",X"C8",X"4F",X"23",X"5E",X"23",X"56",X"EB",X"3E",X"90",X"CD",X"DE",X"3C",X"3E",
		X"01",X"CD",X"F4",X"3C",X"11",X"60",X"00",X"19",X"0D",X"20",X"EF",X"00",X"C9",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"19",X"4E",X"A7",X"C8",X"4F",X"21",X"C1",X"40",X"CD",
		X"6A",X"8C",X"C9",X"3E",X"05",X"CD",X"AB",X"3E",X"3E",X"70",X"CF",X"CD",X"BA",X"2F",X"C9",X"AF",
		X"32",X"9C",X"4E",X"CD",X"41",X"8D",X"CD",X"8B",X"8E",X"32",X"80",X"50",X"CD",X"F6",X"28",X"3E",
		X"11",X"CD",X"AB",X"3E",X"3A",X"70",X"4E",X"21",X"00",X"00",X"22",X"EB",X"90",X"C9",X"FF",X"FF",
		X"21",X"FB",X"4D",X"7E",X"A7",X"C8",X"4F",X"2A",X"17",X"4E",X"11",X"60",X"00",X"ED",X"52",X"22",
		X"17",X"4E",X"0D",X"20",X"F5",X"C9",X"CD",X"09",X"86",X"21",X"19",X"4E",X"34",X"21",X"FB",X"4D",
		X"35",X"CD",X"26",X"8C",X"3A",X"19",X"4E",X"FE",X"07",X"C0",X"3E",X"01",X"32",X"A5",X"4D",X"32",
		X"E2",X"90",X"CD",X"FD",X"8C",X"01",X"06",X"00",X"CD",X"54",X"8C",X"C9",X"FF",X"21",X"00",X"00",
		X"22",X"A7",X"4D",X"22",X"A9",X"4D",X"21",X"E5",X"4D",X"AF",X"06",X"1B",X"CF",X"C9",X"CD",X"FD",
		X"8C",X"CD",X"51",X"8C",X"21",X"04",X"4E",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"C4",X"87",X"22",X"00",X"4D",X"21",X"38",X"2E",X"22",X"0A",X"4D",X"22",X"31",X"4D",X"21",
		X"00",X"FF",X"22",X"14",X"4D",X"22",X"1E",X"4D",X"3E",X"00",X"32",X"28",X"4D",X"32",X"2C",X"4D",
		X"C9",X"3A",X"FB",X"4D",X"A7",X"C8",X"21",X"16",X"4E",X"86",X"77",X"3A",X"FB",X"4D",X"CD",X"C6",
		X"8C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"36",X"A6",X"E5",X"11",X"00",X"04",X"19",X"36",
		X"01",X"E1",X"C9",X"FF",X"FF",X"FF",X"3A",X"FB",X"4D",X"A7",X"28",X"0B",X"21",X"16",X"4E",X"86",
		X"77",X"3A",X"FB",X"4D",X"CD",X"C6",X"8C",X"21",X"16",X"4E",X"CD",X"60",X"8C",X"CD",X"D0",X"A4",
		X"C9",X"CD",X"C0",X"3E",X"21",X"16",X"4E",X"CD",X"60",X"8C",X"CD",X"86",X"8C",X"3E",X"03",X"32",
		X"80",X"50",X"CD",X"DB",X"80",X"CD",X"EE",X"80",X"C9",X"3A",X"FE",X"4D",X"A7",X"28",X"07",X"AF",
		X"32",X"FE",X"4D",X"CD",X"B3",X"8D",X"3A",X"FF",X"4D",X"A7",X"C8",X"AF",X"32",X"FF",X"4D",X"CD",
		X"B3",X"8D",X"C9",X"3A",X"A5",X"4D",X"A7",X"C0",X"21",X"FB",X"4D",X"7E",X"A7",X"C8",X"35",X"CD",
		X"49",X"8C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"9C",X"A6",X"78",X"FE",X"05",
		X"20",X"02",X"3D",X"05",X"32",X"A4",X"4D",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"EA",X"90",X"A7",X"20",X"04",
		X"21",X"3E",X"3D",X"C9",X"21",X"F7",X"8B",X"C9",X"CD",X"A6",X"8E",X"21",X"00",X"90",X"06",X"0F",
		X"AF",X"CF",X"21",X"00",X"00",X"22",X"F0",X"90",X"22",X"F2",X"90",X"C9",X"F5",X"ED",X"57",X"B7",
		X"28",X"04",X"F1",X"C3",X"D4",X"3B",X"F1",X"C3",X"30",X"3D",X"FF",X"CD",X"C2",X"1F",X"3E",X"5C",
		X"32",X"9D",X"41",X"3E",X"01",X"32",X"9D",X"45",X"06",X"17",X"CD",X"5E",X"2C",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"CD",X"51",X"8C",X"3A",X"13",X"4E",X"A7",X"C0",X"CD",X"00",X"81",X"C9",X"FF",X"FF",
		X"06",X"01",X"CD",X"ED",X"23",X"CD",X"D7",X"24",X"CD",X"B3",X"8D",X"AF",X"21",X"E0",X"4D",X"06",
		X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",X"CF",X"CD",X"81",X"8D",X"CD",X"7F",X"0F",X"CD",X"08",
		X"8E",X"CD",X"77",X"25",X"C9",X"06",X"03",X"CD",X"5A",X"2A",X"CD",X"D2",X"8A",X"C3",X"40",X"19",
		X"FE",X"03",X"CA",X"C2",X"8B",X"3E",X"01",X"32",X"E2",X"90",X"C9",X"AF",X"21",X"E0",X"4D",X"06",
		X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",X"CF",X"C9",X"FF",X"3E",X"01",X"32",X"80",X"50",X"3A",
		X"F6",X"4D",X"C9",X"CD",X"C0",X"3E",X"3A",X"1C",X"4E",X"CD",X"19",X"81",X"C9",X"3A",X"E4",X"4D",
		X"FE",X"01",X"CA",X"76",X"01",X"FE",X"02",X"28",X"06",X"CD",X"9E",X"84",X"C3",X"76",X"01",X"CD",
		X"D0",X"8E",X"C3",X"76",X"01",X"AF",X"32",X"E4",X"4D",X"CD",X"CC",X"81",X"CD",X"8B",X"87",X"C9",
		X"2A",X"22",X"4C",X"ED",X"5B",X"2A",X"4C",X"22",X"2A",X"4C",X"ED",X"53",X"22",X"4C",X"CD",X"64",
		X"8F",X"ED",X"5B",X"3A",X"4C",X"22",X"3A",X"4C",X"ED",X"53",X"32",X"4C",X"C9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"48",X"4D",X"7E",X"8F",X"77",X"C9",X"21",X"4C",
		X"3E",X"9E",X"21",X"11",X"42",X"CD",X"DE",X"3C",X"3E",X"01",X"CD",X"F4",X"3C",X"C9",X"FF",X"FF",
		X"CD",X"9E",X"85",X"CD",X"10",X"81",X"C9",X"CD",X"66",X"8D",X"CD",X"A6",X"0A",X"3A",X"09",X"4E",
		X"EE",X"01",X"32",X"09",X"4E",X"C3",X"6C",X"09",X"3A",X"01",X"90",X"A7",X"28",X"07",X"78",X"FE",
		X"04",X"C8",X"FE",X"03",X"C8",X"3A",X"02",X"90",X"A7",X"38",X"07",X"78",X"FE",X"02",X"C8",X"FE",
		X"01",X"C8",X"CD",X"CF",X"88",X"C9",X"3A",X"03",X"90",X"A7",X"28",X"07",X"78",X"FE",X"04",X"C8",
		X"FE",X"03",X"C8",X"3A",X"04",X"90",X"A7",X"28",X"07",X"78",X"FE",X"02",X"C8",X"FE",X"01",X"C8",
		X"CD",X"CF",X"88",X"C9",X"21",X"32",X"4C",X"34",X"2A",X"32",X"4C",X"C9",X"CA",X"B6",X"8B",X"05",
		X"2A",X"D2",X"4D",X"3E",X"10",X"95",X"ED",X"5B",X"08",X"4D",X"A7",X"ED",X"52",X"CA",X"B6",X"8B",
		X"C3",X"08",X"3B",X"3E",X"01",X"32",X"A8",X"4D",X"32",X"AD",X"4D",X"C9",X"CD",X"70",X"84",X"0E",
		X"03",X"3E",X"76",X"21",X"BC",X"41",X"CD",X"DE",X"3C",X"F5",X"3E",X"01",X"CD",X"F4",X"3C",X"F1",
		X"06",X"04",X"80",X"11",X"40",X"00",X"19",X"0D",X"20",X"EC",X"CD",X"2B",X"8E",X"C9",X"00",X"00",
		X"C4",X"40",X"16",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"6C",X"08",X"07",X"00",X"00",X"06",
		X"05",X"00",X"04",X"03",X"02",X"01",X"FE",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"6D",X"1F",X"1E",
		X"1D",X"1C",X"00",X"00",X"00",X"1B",X"00",X"1A",X"19",X"18",X"17",X"FE",X"6B",X"6A",X"69",X"68",
		X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"00",X"00",X"60",X"3F",X"3E",X"3D",X"3C",X"2F",X"2E",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"04",X"02",X"01",X"03",X"02",X"04",X"02",X"03",X"04",X"01",X"01",X"02",X"04",X"03",
		X"02",X"03",X"01",X"04",X"03",X"02",X"04",X"01",X"01",X"01",X"03",X"04",X"02",X"01",X"04",X"03",
		X"03",X"02",X"01",X"04",X"04",X"02",X"03",X"01",X"02",X"01",X"03",X"04",X"03",X"01",X"04",X"02",
		X"04",X"02",X"01",X"03",X"03",X"01",X"02",X"04",X"04",X"01",X"03",X"02",X"04",X"01",X"02",X"03",
		X"00",X"04",X"08",X"0C",X"10",X"14",X"18",X"1C",X"20",X"24",X"28",X"2C",X"30",X"34",X"38",X"3C",
		X"F5",X"E5",X"D5",X"3A",X"C0",X"50",X"E6",X"0F",X"5F",X"16",X"00",X"21",X"40",X"80",X"19",X"5E",
		X"21",X"00",X"80",X"19",X"11",X"E0",X"4D",X"01",X"04",X"00",X"ED",X"B0",X"D1",X"E1",X"F1",X"C9",
		X"F5",X"AF",X"32",X"80",X"50",X"00",X"00",X"00",X"F1",X"C9",X"CD",X"0F",X"20",X"FE",X"FC",X"28",
		X"02",X"FE",X"FD",X"CA",X"40",X"19",X"FE",X"70",X"C3",X"F0",X"88",X"7D",X"21",X"E0",X"4D",X"FE",
		X"EB",X"28",X"14",X"FE",X"90",X"20",X"03",X"23",X"18",X"0D",X"FE",X"F4",X"20",X"04",X"23",X"23",
		X"18",X"05",X"FE",X"70",X"23",X"23",X"23",X"7E",X"32",X"E4",X"4D",X"3E",X"72",X"CD",X"9E",X"3E",
		X"3E",X"11",X"CD",X"AB",X"3E",X"C3",X"75",X"8E",X"FF",X"FF",X"FF",X"3A",X"E6",X"4D",X"A7",X"C0",
		X"3E",X"01",X"32",X"E6",X"4D",X"CD",X"3D",X"81",X"CD",X"2D",X"83",X"C9",X"3E",X"01",X"06",X"03",
		X"11",X"20",X"00",X"C5",X"D5",X"E5",X"CF",X"E1",X"D1",X"C1",X"C9",X"21",X"CD",X"45",X"CD",X"CC",
		X"80",X"19",X"CD",X"CC",X"80",X"19",X"CD",X"CC",X"80",X"19",X"CD",X"CC",X"80",X"C9",X"01",X"FD",
		X"80",X"21",X"D0",X"41",X"CD",X"72",X"81",X"3E",X"DA",X"32",X"30",X"42",X"C9",X"DA",X"DA",X"DA",
		X"CD",X"69",X"8B",X"CD",X"77",X"8D",X"CD",X"DB",X"80",X"CD",X"EE",X"80",X"C9",X"00",X"00",X"00",
		X"3A",X"1C",X"4E",X"C6",X"99",X"27",X"CD",X"A8",X"85",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"C6",
		X"30",X"32",X"F2",X"41",X"3A",X"1C",X"4E",X"E6",X"0F",X"C6",X"30",X"32",X"D2",X"41",X"3E",X"0F",
		X"32",X"F2",X"45",X"32",X"D2",X"45",X"CD",X"B2",X"82",X"C9",X"F0",X"72",X"F1",X"3E",X"11",X"CD",
		X"99",X"0F",X"01",X"3A",X"81",X"21",X"84",X"40",X"CD",X"72",X"81",X"21",X"64",X"41",X"CD",X"72",
		X"81",X"21",X"44",X"42",X"CD",X"72",X"81",X"21",X"24",X"43",X"CD",X"72",X"81",X"C9",X"3E",X"17",
		X"CD",X"99",X"0F",X"01",X"ED",X"0F",X"CD",X"45",X"81",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"C5",X"00",X"11",X"20",X"00",X"0A",X"77",X"19",X"03",X"0A",X"77",X"19",X"03",X"0A",
		X"77",X"C1",X"C9",X"3A",X"FA",X"4D",X"A7",X"C0",X"3A",X"E6",X"4D",X"A7",X"C0",X"3E",X"01",X"32",
		X"E6",X"4D",X"CD",X"3D",X"81",X"CD",X"2D",X"83",X"21",X"9C",X"4E",X"36",X"10",X"C9",X"21",X"BC",
		X"4E",X"36",X"02",X"21",X"04",X"4E",X"C9",X"21",X"90",X"4C",X"3A",X"8A",X"4C",X"4F",X"06",X"10",
		X"7E",X"A7",X"28",X"2F",X"E6",X"C0",X"07",X"07",X"B9",X"30",X"28",X"35",X"7E",X"E6",X"3F",X"20",
		X"22",X"77",X"C5",X"E5",X"2C",X"7E",X"2C",X"46",X"21",X"E1",X"81",X"E5",X"E7",X"94",X"08",X"A3",
		X"06",X"8E",X"05",X"42",X"12",X"00",X"10",X"0B",X"10",X"63",X"02",X"2B",X"21",X"F0",X"21",X"B9",
		X"22",X"E1",X"C1",X"2C",X"2C",X"2C",X"10",X"C8",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"3A",X"ED",X"4D",X"A7",X"20",X"09",X"3E",X"01",X"32",X"ED",X"4D",X"CD",X"E9",
		X"0F",X"C9",X"3A",X"EF",X"4D",X"A7",X"20",X"04",X"CD",X"79",X"3F",X"C9",X"C3",X"61",X"84",X"00",
		X"21",X"00",X"40",X"CF",X"06",X"3F",X"21",X"C0",X"43",X"CF",X"3A",X"EE",X"4D",X"A7",X"C0",X"3E",
		X"01",X"32",X"E8",X"4D",X"CD",X"82",X"3C",X"C9",X"3A",X"E8",X"4D",X"A7",X"C0",X"3A",X"09",X"4E",
		X"C3",X"47",X"03",X"CD",X"3E",X"75",X"21",X"37",X"43",X"11",X"20",X"00",X"77",X"3D",X"19",X"77",
		X"3E",X"05",X"32",X"37",X"47",X"32",X"57",X"47",X"CD",X"8A",X"05",X"C9",X"1F",X"C9",X"AF",X"32",
		X"B1",X"4D",X"C9",X"F1",X"02",X"F2",X"03",X"F3",X"0F",X"70",X"F4",X"02",X"8D",X"F4",X"02",X"88",
		X"F4",X"02",X"8A",X"70",X"F4",X"01",X"6C",X"F4",X"02",X"8A",X"F4",X"01",X"6A",X"F4",X"02",X"88",
		X"70",X"F4",X"02",X"8D",X"F4",X"02",X"88",X"F4",X"02",X"8A",X"70",X"F4",X"01",X"6C",X"F4",X"02",
		X"8A",X"F4",X"01",X"6A",X"F4",X"02",X"88",X"70",X"F0",X"6A",X"82",X"FF",X"21",X"BC",X"4E",X"CB",
		X"AE",X"3E",X"01",X"32",X"F5",X"90",X"C9",X"3E",X"01",X"32",X"F4",X"90",X"CD",X"9C",X"82",X"CB",
		X"F6",X"C9",X"3A",X"EA",X"90",X"A7",X"C0",X"CD",X"00",X"8F",X"C9",X"3E",X"01",X"32",X"80",X"50",
		X"C9",X"3E",X"00",X"32",X"80",X"50",X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"28",X"10",X"AF",X"32",
		X"80",X"50",X"CD",X"51",X"8C",X"CD",X"00",X"81",X"3E",X"02",X"32",X"80",X"50",X"C9",X"3A",X"1C",
		X"4E",X"A7",X"20",X"10",X"CD",X"C0",X"8C",X"3A",X"FB",X"4D",X"21",X"16",X"4E",X"86",X"77",X"3E",
		X"40",X"32",X"1C",X"4E",X"AF",X"21",X"E0",X"4D",X"06",X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",
		X"CF",X"CD",X"00",X"81",X"CD",X"35",X"A4",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"21",
		X"00",X"00",X"22",X"FC",X"4D",X"22",X"FE",X"4D",X"C9",X"CD",X"7C",X"0E",X"3E",X"20",X"32",X"04",
		X"4E",X"C9",X"CD",X"6C",X"0E",X"CD",X"B0",X"0E",X"CD",X"C1",X"2C",X"C9",X"FF",X"06",X"16",X"CD",
		X"5E",X"2C",X"C9",X"FF",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"08",X"DD",X"21",X"E9",X"4D",X"C9",
		X"DD",X"21",X"39",X"4D",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"06",X"3A",X"AF",X"4D",X"C3",
		X"4C",X"3D",X"3A",X"AC",X"4D",X"A7",X"28",X"06",X"3A",X"AF",X"4D",X"C3",X"4C",X"3D",X"3A",X"F9",
		X"4D",X"A7",X"C2",X"83",X"83",X"3A",X"16",X"4E",X"A7",X"CA",X"4C",X"83",X"2A",X"31",X"4D",X"11",
		X"22",X"23",X"A7",X"ED",X"52",X"C2",X"4C",X"83",X"3E",X"08",X"32",X"F9",X"4D",X"C3",X"4C",X"83",
		X"00",X"00",X"00",X"2A",X"31",X"4D",X"11",X"3A",X"2D",X"A7",X"ED",X"52",X"C2",X"4C",X"83",X"AF",
		X"32",X"F9",X"4D",X"C3",X"45",X"83",X"00",X"00",X"00",X"3A",X"E4",X"4D",X"FE",X"01",X"C2",X"02",
		X"3E",X"3E",X"01",X"32",X"A7",X"4D",X"C3",X"63",X"17",X"2A",X"39",X"4D",X"7D",X"06",X"23",X"90",
		X"3A",X"39",X"4D",X"D8",X"06",X"25",X"90",X"D8",X"CD",X"D6",X"A0",X"C9",X"FF",X"FF",X"CD",X"FB",
		X"83",X"21",X"00",X"00",X"28",X"03",X"22",X"FC",X"4D",X"22",X"FE",X"4D",X"C9",X"00",X"00",X"00",
		X"00",X"E5",X"D5",X"11",X"20",X"00",X"77",X"3C",X"19",X"77",X"3C",X"3C",X"23",X"77",X"3D",X"ED",
		X"52",X"77",X"D1",X"E1",X"C9",X"CD",X"17",X"2D",X"3A",X"00",X"4E",X"FE",X"03",X"D0",X"CD",X"F3",
		X"2C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"E4",X"4D",X"FE",X"01",
		X"C9",X"FD",X"21",X"0A",X"4D",X"CD",X"FB",X"83",X"28",X"09",X"DD",X"21",X"E9",X"4D",X"CD",X"FA",
		X"09",X"18",X"03",X"CD",X"A9",X"31",X"30",X"0E",X"3A",X"B1",X"4D",X"A7",X"C0",X"3E",X"01",X"32",
		X"B1",X"4D",X"CD",X"07",X"1F",X"C9",X"AF",X"32",X"B1",X"4D",X"C9",X"F5",X"E5",X"D5",X"11",X"00",
		X"04",X"3E",X"11",X"19",X"77",X"D1",X"E1",X"F1",X"77",X"C9",X"D5",X"E5",X"06",X"20",X"4F",X"CD",
		X"2B",X"84",X"F5",X"E5",X"11",X"E0",X"83",X"7D",X"E6",X"1F",X"87",X"26",X"00",X"6F",X"19",X"D1",
		X"A7",X"ED",X"52",X"F1",X"EE",X"01",X"CD",X"2B",X"84",X"EB",X"23",X"79",X"10",X"E1",X"E1",X"D1",
		X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"C2",X"2A",X"82",X"3E",X"40",X"06",X"3F",X"C3",X"20",X"82",
		X"2A",X"B0",X"8F",X"22",X"86",X"4D",X"11",X"B2",X"8F",X"01",X"20",X"00",X"1A",X"FE",X"FF",X"C8",
		X"FE",X"FE",X"20",X"0A",X"2A",X"86",X"4D",X"23",X"22",X"86",X"4D",X"13",X"18",X"EE",X"77",X"E5",
		X"C5",X"01",X"00",X"04",X"09",X"3E",X"01",X"77",X"C1",X"E1",X"09",X"13",X"18",X"DE",X"2A",X"24",
		X"4C",X"ED",X"5B",X"26",X"4C",X"ED",X"4B",X"28",X"4C",X"22",X"26",X"4C",X"ED",X"53",X"28",X"4C",
		X"2A",X"2A",X"4C",X"ED",X"43",X"2A",X"4C",X"22",X"24",X"4C",X"2A",X"34",X"4C",X"ED",X"5B",X"36",
		X"4C",X"ED",X"4B",X"38",X"4C",X"22",X"36",X"4C",X"ED",X"53",X"38",X"4C",X"2A",X"3A",X"4C",X"ED",
		X"43",X"3A",X"4C",X"22",X"34",X"4C",X"C9",X"21",X"83",X"E3",X"22",X"02",X"4D",X"21",X"83",X"D1",
		X"22",X"04",X"4D",X"21",X"83",X"BF",X"22",X"06",X"4D",X"CD",X"99",X"14",X"C9",X"21",X"97",X"D1",
		X"22",X"00",X"4D",X"CD",X"99",X"14",X"C9",X"3E",X"94",X"21",X"34",X"43",X"77",X"E5",X"23",X"3C",
		X"77",X"23",X"3C",X"77",X"E1",X"11",X"20",X"00",X"19",X"3C",X"77",X"23",X"3C",X"77",X"23",X"3C",
		X"77",X"3E",X"01",X"21",X"34",X"47",X"11",X"20",X"00",X"01",X"00",X"03",X"E5",X"C5",X"CF",X"C1",
		X"E1",X"19",X"CF",X"C9",X"3E",X"01",X"CD",X"74",X"0F",X"C9",X"01",X"5A",X"85",X"CD",X"72",X"81",
		X"C9",X"E5",X"CD",X"2A",X"85",X"E1",X"11",X"00",X"04",X"19",X"CD",X"24",X"85",X"C9",X"21",X"50",
		X"40",X"CD",X"31",X"85",X"C9",X"21",X"53",X"40",X"CD",X"31",X"85",X"C9",X"21",X"55",X"40",X"CD",
		X"31",X"85",X"C9",X"21",X"57",X"40",X"CD",X"31",X"85",X"C9",X"53",X"54",X"50",X"AF",X"32",X"FB",
		X"4D",X"21",X"00",X"00",X"22",X"A4",X"4D",X"21",X"31",X"93",X"22",X"08",X"4D",X"CD",X"99",X"14",
		X"06",X"01",X"CD",X"ED",X"23",X"CD",X"B3",X"85",X"CD",X"8A",X"05",X"C9",X"21",X"FB",X"4D",X"19",
		X"D5",X"E5",X"11",X"A7",X"4D",X"A7",X"ED",X"52",X"E1",X"D1",X"06",X"02",X"28",X"0A",X"06",X"00",
		X"7E",X"A7",X"28",X"07",X"06",X"01",X"AF",X"77",X"CD",X"CD",X"0F",X"CD",X"10",X"81",X"CD",X"5A",
		X"2A",X"CD",X"12",X"86",X"00",X"E6",X"C9",X"C9",X"32",X"1C",X"4E",X"A7",X"C0",X"3E",X"01",X"32",
		X"DF",X"90",X"C9",X"CD",X"70",X"84",X"CD",X"38",X"8E",X"C9",X"FF",X"FF",X"21",X"00",X"00",X"22",
		X"08",X"4D",X"22",X"02",X"4D",X"22",X"04",X"4D",X"22",X"06",X"4D",X"22",X"00",X"4D",X"22",X"F0",
		X"90",X"22",X"F2",X"90",X"22",X"D2",X"4D",X"22",X"E4",X"4D",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",
		X"20",X"04",X"CD",X"56",X"89",X"C9",X"FE",X"02",X"20",X"07",X"CD",X"70",X"8B",X"CD",X"49",X"3D",
		X"C9",X"06",X"04",X"ED",X"5B",X"39",X"4D",X"CD",X"23",X"17",X"CD",X"49",X"3D",X"C9",X"21",X"BC",
		X"4E",X"CB",X"DE",X"CD",X"9C",X"82",X"C9",X"FF",X"FF",X"21",X"BC",X"4E",X"CB",X"D6",X"CD",X"9C",
		X"82",X"C9",X"21",X"BC",X"4E",X"36",X"10",X"CD",X"9C",X"82",X"CD",X"17",X"2D",X"C9",X"FF",X"FF",
		X"CD",X"FB",X"83",X"28",X"07",X"DD",X"21",X"01",X"33",X"C3",X"D6",X"10",X"EF",X"04",X"01",X"AF",
		X"32",X"AC",X"4D",X"32",X"A7",X"4D",X"32",X"F0",X"90",X"C3",X"01",X"11",X"21",X"F0",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"4F",X"1B",X"C3",X"C3",X"10",X"21",X"F1",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"C7",X"1B",X"C3",X"1B",X"11",X"21",X"F2",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"3F",X"1C",X"C3",X"5F",X"11",X"21",X"F3",X"90",X"7E",
		X"FE",X"F0",X"28",X"02",X"34",X"C9",X"CD",X"B7",X"1C",X"C3",X"CC",X"11",X"3A",X"E4",X"4D",X"32",
		X"FF",X"90",X"C9",X"3A",X"00",X"4E",X"FE",X"03",X"D0",X"3E",X"02",X"32",X"9C",X"4E",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"21",X"06",X"4C",X"06",X"04",X"1A",X"77",X"23",X"23",X"13",X"05",X"20",
		X"F8",X"C9",X"21",X"07",X"4C",X"3E",X"09",X"06",X"04",X"77",X"23",X"23",X"05",X"20",X"FA",X"C9",
		X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"C9",X"CD",X"3F",X"88",X"11",X"61",X"12",X"A7",
		X"C8",X"11",X"65",X"12",X"C9",X"CD",X"33",X"88",X"11",X"69",X"12",X"A7",X"C8",X"11",X"6D",X"12",
		X"C9",X"CD",X"57",X"88",X"11",X"71",X"12",X"A7",X"C8",X"11",X"75",X"12",X"C9",X"CD",X"4B",X"88",
		X"11",X"79",X"12",X"A7",X"C8",X"11",X"7D",X"12",X"C9",X"CD",X"B0",X"86",X"20",X"22",X"3A",X"30",
		X"4D",X"FE",X"00",X"20",X"04",X"CD",X"C5",X"86",X"C9",X"FE",X"01",X"20",X"04",X"CD",X"B9",X"86",
		X"C9",X"FE",X"02",X"20",X"04",X"CD",X"B9",X"86",X"C9",X"FE",X"03",X"C0",X"CD",X"C5",X"86",X"C9",
		X"3A",X"30",X"4D",X"FE",X"00",X"20",X"04",X"CD",X"DD",X"86",X"C9",X"FE",X"01",X"20",X"04",X"CD",
		X"D1",X"86",X"C9",X"FE",X"02",X"20",X"04",X"CD",X"D1",X"86",X"C9",X"FE",X"03",X"C0",X"CD",X"DD",
		X"86",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"04",X"CD",X"9C",X"16",X"C9",X"CD",X"E9",X"86",
		X"CD",X"94",X"86",X"CD",X"A2",X"86",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"04",X"CD",X"AA",
		X"16",X"C9",X"CD",X"E9",X"86",X"CD",X"94",X"86",X"CD",X"A2",X"86",X"C9",X"21",X"02",X"4C",X"CD",
		X"4E",X"15",X"CD",X"32",X"87",X"CD",X"47",X"87",X"C9",X"21",X"00",X"00",X"22",X"01",X"90",X"22",
		X"03",X"90",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"28",X"08",X"FE",X"02",X"28",X"04",X"CD",X"09",
		X"3D",X"C9",X"3A",X"FD",X"4D",X"A7",X"C8",X"CD",X"09",X"3D",X"C9",X"3E",X"40",X"06",X"0C",X"21",
		X"45",X"41",X"CD",X"76",X"0F",X"C9",X"00",X"DD",X"21",X"26",X"4D",X"CD",X"0F",X"20",X"21",X"00",
		X"90",X"FE",X"FC",X"28",X"0D",X"FE",X"FD",X"28",X"09",X"E6",X"C0",X"D6",X"C0",X"20",X"03",X"36",
		X"01",X"C9",X"36",X"00",X"C9",X"0D",X"0C",X"0B",X"0A",X"09",X"6C",X"08",X"07",X"00",X"00",X"06",
		X"2A",X"39",X"4D",X"7D",X"06",X"02",X"80",X"32",X"D2",X"4D",X"7C",X"32",X"D3",X"4D",X"C9",X"1E",
		X"3A",X"3C",X"4D",X"FE",X"00",X"20",X"12",X"FD",X"21",X"35",X"4D",X"CD",X"97",X"87",X"7E",X"A7",
		X"C0",X"FD",X"21",X"37",X"4D",X"CD",X"97",X"87",X"C9",X"FE",X"01",X"20",X"15",X"CD",X"C0",X"87",
		X"FD",X"21",X"D2",X"4D",X"CD",X"97",X"87",X"7E",X"A7",X"C0",X"FD",X"21",X"37",X"4D",X"CD",X"97",
		X"87",X"C9",X"FE",X"02",X"20",X"04",X"CD",X"ED",X"87",X"C9",X"FE",X"03",X"C0",X"CD",X"D7",X"87",
		X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"08",X"CD",X"D0",X"87",X"3A",X"00",X"90",X"A7",X"C0",
		X"FD",X"21",X"39",X"4D",X"C3",X"7A",X"80",X"AF",X"21",X"00",X"90",X"01",X"FF",X"03",X"CF",X"C3",
		X"3E",X"A7",X"00",X"CD",X"69",X"87",X"3E",X"01",X"32",X"01",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",
		X"69",X"87",X"3E",X"01",X"32",X"02",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",X"69",X"87",X"3E",X"01",
		X"32",X"03",X"90",X"3A",X"C0",X"4D",X"C9",X"CD",X"69",X"87",X"3E",X"01",X"32",X"04",X"90",X"3A",
		X"C0",X"4D",X"C9",X"06",X"04",X"2A",X"37",X"4D",X"A7",X"ED",X"52",X"28",X"1C",X"05",X"2A",X"35",
		X"4D",X"A7",X"ED",X"52",X"28",X"13",X"05",X"2A",X"39",X"4D",X"A7",X"ED",X"52",X"28",X"0A",X"05",
		X"2A",X"D2",X"4D",X"A7",X"ED",X"52",X"28",X"01",X"05",X"78",X"C9",X"3A",X"FD",X"4D",X"A7",X"3E",
		X"01",X"28",X"03",X"32",X"FB",X"4D",X"32",X"FF",X"90",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"ED",X"5B",X"33",X"4D",X"CD",X"63",X"88",X"32",X"06",X"90",X"A7",X"C8",X"3E",X"01",X"32",X"A8",
		X"4D",X"3E",X"02",X"32",X"A4",X"4D",X"C9",X"ED",X"5B",X"31",X"4D",X"CD",X"63",X"88",X"32",X"05",
		X"90",X"A7",X"C8",X"3E",X"01",X"32",X"A7",X"4D",X"32",X"A4",X"4D",X"C9",X"00",X"00",X"00",X"3A",
		X"05",X"90",X"A7",X"28",X"0B",X"AF",X"32",X"A7",X"4D",X"32",X"05",X"90",X"32",X"A4",X"4D",X"C9",
		X"3A",X"06",X"90",X"A7",X"C8",X"AF",X"32",X"A8",X"4D",X"32",X"06",X"90",X"32",X"A4",X"4D",X"C9",
		X"CA",X"8B",X"80",X"FE",X"90",X"CA",X"F5",X"18",X"FE",X"92",X"CA",X"F5",X"18",X"C3",X"EF",X"18",
		X"A7",X"C8",X"47",X"CD",X"B0",X"86",X"20",X"04",X"CD",X"28",X"8F",X"C9",X"CD",X"46",X"8F",X"C9",
		X"31",X"C0",X"4F",X"AF",X"01",X"04",X"00",X"21",X"00",X"90",X"CF",X"0D",X"20",X"FC",X"C3",X"3E",
		X"A7",X"00",X"00",X"00",X"C8",X"78",X"FE",X"02",X"C8",X"FE",X"01",X"C8",X"3E",X"01",X"32",X"A4",
		X"4D",X"CD",X"CF",X"88",X"C9",X"D6",X"C0",X"28",X"0A",X"7E",X"FE",X"90",X"28",X"05",X"FE",X"92",
		X"C2",X"9F",X"29",X"11",X"00",X"04",X"19",X"7E",X"FE",X"16",X"CA",X"0B",X"8B",X"FE",X"17",X"CA",
		X"9F",X"29",X"C3",X"C6",X"29",X"FF",X"3A",X"AC",X"4D",X"A7",X"C0",X"00",X"00",X"CD",X"B7",X"88",
		X"3A",X"05",X"90",X"CD",X"00",X"89",X"A7",X"28",X"09",X"AF",X"32",X"08",X"90",X"06",X"02",X"CD",
		X"9B",X"85",X"CD",X"49",X"3D",X"3A",X"AD",X"4D",X"A7",X"C0",X"00",X"00",X"CD",X"A0",X"88",X"3A",
		X"06",X"90",X"CD",X"00",X"89",X"A7",X"20",X"06",X"CD",X"49",X"3D",X"C9",X"00",X"00",X"3A",X"A4",
		X"4D",X"CD",X"6C",X"17",X"AF",X"32",X"FD",X"4D",X"CD",X"49",X"3D",X"C9",X"00",X"00",X"00",X"00",
		X"21",X"02",X"4C",X"CD",X"4E",X"15",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"07",X"CD",X"32",X"87",
		X"CD",X"47",X"87",X"C9",X"FE",X"02",X"C0",X"CD",X"E0",X"89",X"C9",X"00",X"00",X"00",X"00",X"00",
		X"5E",X"23",X"56",X"23",X"4E",X"23",X"46",X"C9",X"CD",X"C0",X"89",X"ED",X"53",X"02",X"4C",X"ED",
		X"43",X"06",X"4C",X"23",X"CD",X"C0",X"89",X"ED",X"53",X"08",X"4C",X"ED",X"43",X"0C",X"4C",X"C9",
		X"3A",X"E4",X"4D",X"FE",X"02",X"C0",X"CD",X"B0",X"86",X"20",X"10",X"3A",X"C0",X"4D",X"21",X"10",
		X"8A",X"A7",X"20",X"03",X"21",X"18",X"8A",X"CD",X"C8",X"89",X"C9",X"3A",X"C0",X"4D",X"21",X"20",
		X"8A",X"A7",X"20",X"03",X"21",X"28",X"8A",X"CD",X"C8",X"89",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"68",X"01",X"60",X"01",X"64",X"01",X"6C",X"01",X"78",X"01",X"70",X"01",X"74",X"01",X"7C",X"01",
		X"6B",X"01",X"63",X"01",X"67",X"01",X"6F",X"01",X"7B",X"01",X"73",X"01",X"77",X"01",X"7F",X"01",
		X"3E",X"FD",X"21",X"85",X"40",X"06",X"15",X"CF",X"21",X"B9",X"40",X"11",X"20",X"00",X"06",X"18",
		X"77",X"19",X"05",X"20",X"FB",X"21",X"8A",X"42",X"06",X"0A",X"CF",X"00",X"00",X"00",X"00",X"21",
		X"CA",X"41",X"06",X"06",X"77",X"19",X"05",X"20",X"FB",X"21",X"AA",X"41",X"77",X"23",X"77",X"21",
		X"73",X"42",X"77",X"C3",X"50",X"8B",X"AF",X"06",X"5F",X"21",X"8C",X"4E",X"CF",X"C9",X"FF",X"FF",
		X"3E",X"40",X"21",X"A5",X"40",X"06",X"14",X"CF",X"21",X"A9",X"42",X"06",X"0B",X"CF",X"21",X"D8",
		X"40",X"06",X"17",X"77",X"19",X"05",X"20",X"FB",X"21",X"A9",X"41",X"06",X"08",X"77",X"19",X"05",
		X"20",X"FB",X"21",X"89",X"41",X"77",X"23",X"77",X"21",X"6F",X"40",X"77",X"23",X"77",X"C9",X"FF",
		X"84",X"44",X"85",X"44",X"88",X"44",X"8E",X"44",X"91",X"44",X"97",X"44",X"39",X"45",X"99",X"45",
		X"79",X"46",X"D9",X"46",X"99",X"47",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"06",X"0B",X"11",X"A0",X"8A",X"1A",X"6F",X"13",X"1A",X"67",X"3E",X"16",X"77",X"13",X"05",X"20",
		X"F4",X"C9",X"3A",X"E4",X"4D",X"FE",X"01",X"20",X"07",X"CD",X"00",X"81",X"CD",X"3D",X"25",X"C9",
		X"FE",X"02",X"C0",X"CD",X"00",X"81",X"CD",X"30",X"8A",X"CD",X"70",X"8A",X"CD",X"C0",X"8A",X"CD",
		X"20",X"8D",X"C9",X"FE",X"90",X"CA",X"23",X"19",X"FE",X"92",X"CA",X"23",X"19",X"E6",X"C0",X"D6",
		X"C0",X"CA",X"23",X"19",X"C3",X"50",X"19",X"FF",X"FF",X"FF",X"FF",X"DD",X"E5",X"FD",X"E5",X"00",
		X"00",X"00",X"00",X"FD",X"21",X"0C",X"4D",X"CD",X"0F",X"20",X"19",X"7E",X"FD",X"E1",X"DD",X"E1",
		X"FE",X"16",X"CA",X"9F",X"29",X"C3",X"C6",X"29",X"3A",X"E4",X"4D",X"21",X"00",X"00",X"FE",X"02",
		X"28",X"07",X"FE",X"01",X"C0",X"22",X"FE",X"4D",X"C9",X"22",X"FE",X"4D",X"AF",X"32",X"FC",X"4D",
		X"C9",X"BC",X"02",X"5C",X"40",X"53",X"45",X"47",X"41",X"40",X"31",X"39",X"38",X"32",X"2F",X"81",
		X"21",X"D2",X"D2",X"22",X"4F",X"40",X"21",X"FC",X"FC",X"22",X"4F",X"43",X"22",X"6F",X"43",X"22",
		X"8F",X"43",X"21",X"D3",X"D3",X"22",X"AF",X"43",X"C9",X"CD",X"A3",X"8E",X"CD",X"7F",X"0F",X"C9",
		X"06",X"05",X"ED",X"5B",X"39",X"4D",X"3A",X"AF",X"4D",X"A7",X"20",X"09",X"2A",X"37",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AE",X"4D",X"A7",X"20",X"09",X"2A",X"35",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AD",X"4D",X"A7",X"20",X"09",X"2A",X"33",X"4D",X"A7",
		X"ED",X"52",X"CA",X"B6",X"8B",X"05",X"3A",X"AC",X"4D",X"A7",X"20",X"09",X"2A",X"31",X"4D",X"A7",
		X"ED",X"52",X"C3",X"6C",X"8F",X"05",X"CD",X"CD",X"8D",X"00",X"32",X"A5",X"4D",X"A7",X"C8",X"C3",
		X"80",X"8E",X"CD",X"83",X"8F",X"AF",X"32",X"A5",X"4D",X"3A",X"FD",X"4D",X"A7",X"06",X"00",X"28",
		X"09",X"AF",X"32",X"FD",X"4D",X"CD",X"CD",X"0F",X"06",X"01",X"CD",X"10",X"8F",X"C9",X"21",X"02",
		X"4C",X"11",X"F0",X"90",X"06",X"04",X"1A",X"A7",X"28",X"06",X"FE",X"F0",X"20",X"02",X"36",X"FC",
		X"23",X"23",X"13",X"05",X"20",X"F0",X"C9",X"00",X"DD",X"40",X"07",X"C1",X"40",X"40",X"FF",X"FF",
		X"2A",X"17",X"4E",X"3E",X"40",X"CD",X"F4",X"3C",X"11",X"60",X"00",X"19",X"22",X"17",X"4E",X"C9",
		X"2A",X"17",X"4E",X"11",X"60",X"00",X"ED",X"52",X"22",X"17",X"4E",X"3E",X"90",X"CD",X"DE",X"3C",
		X"3E",X"01",X"CD",X"F4",X"3C",X"C9",X"2A",X"1A",X"4E",X"CD",X"1B",X"8C",X"11",X"60",X"00",X"19",
		X"22",X"1A",X"4E",X"C9",X"2A",X"1A",X"4E",X"11",X"60",X"00",X"ED",X"52",X"3E",X"40",X"CD",X"F4",
		X"3C",X"22",X"1A",X"4E",X"C9",X"21",X"FB",X"4D",X"35",X"21",X"16",X"4E",X"34",X"CD",X"10",X"8C",
		X"C9",X"01",X"0B",X"00",X"CD",X"FA",X"8D",X"11",X"16",X"4E",X"ED",X"B0",X"C9",X"00",X"00",X"00",
		X"00",X"7E",X"A7",X"C8",X"4F",X"23",X"5E",X"23",X"56",X"EB",X"3E",X"90",X"CD",X"DE",X"3C",X"3E",
		X"01",X"CD",X"F4",X"3C",X"11",X"60",X"00",X"19",X"0D",X"20",X"EF",X"00",X"C9",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3A",X"19",X"4E",X"A7",X"C8",X"4F",X"21",X"C1",X"40",X"CD",
		X"6A",X"8C",X"C9",X"3E",X"05",X"CD",X"AB",X"3E",X"3E",X"70",X"CF",X"CD",X"BA",X"2F",X"C9",X"AF",
		X"32",X"9C",X"4E",X"CD",X"41",X"8D",X"CD",X"8B",X"8E",X"32",X"80",X"50",X"CD",X"F6",X"28",X"3E",
		X"11",X"CD",X"AB",X"3E",X"3A",X"70",X"4E",X"21",X"00",X"00",X"22",X"EB",X"90",X"C9",X"FF",X"FF",
		X"21",X"FB",X"4D",X"7E",X"A7",X"C8",X"4F",X"2A",X"17",X"4E",X"11",X"60",X"00",X"ED",X"52",X"22",
		X"17",X"4E",X"0D",X"20",X"F5",X"C9",X"CD",X"09",X"86",X"21",X"19",X"4E",X"34",X"21",X"FB",X"4D",
		X"35",X"CD",X"26",X"8C",X"3A",X"19",X"4E",X"FE",X"07",X"C0",X"3E",X"01",X"32",X"A5",X"4D",X"32",
		X"E2",X"90",X"CD",X"FD",X"8C",X"01",X"06",X"00",X"CD",X"54",X"8C",X"C9",X"FF",X"21",X"00",X"00",
		X"22",X"A7",X"4D",X"22",X"A9",X"4D",X"21",X"E5",X"4D",X"AF",X"06",X"1B",X"CF",X"C9",X"CD",X"FD",
		X"8C",X"CD",X"51",X"8C",X"21",X"04",X"4E",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"C4",X"87",X"22",X"00",X"4D",X"21",X"38",X"2E",X"22",X"0A",X"4D",X"22",X"31",X"4D",X"21",
		X"00",X"FF",X"22",X"14",X"4D",X"22",X"1E",X"4D",X"3E",X"00",X"32",X"28",X"4D",X"32",X"2C",X"4D",
		X"C9",X"3A",X"FB",X"4D",X"A7",X"C8",X"21",X"16",X"4E",X"86",X"77",X"3A",X"FB",X"4D",X"CD",X"C6",
		X"8C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"36",X"A6",X"E5",X"11",X"00",X"04",X"19",X"36",
		X"01",X"E1",X"C9",X"FF",X"FF",X"FF",X"3A",X"FB",X"4D",X"A7",X"28",X"0B",X"21",X"16",X"4E",X"86",
		X"77",X"3A",X"FB",X"4D",X"CD",X"C6",X"8C",X"21",X"16",X"4E",X"CD",X"60",X"8C",X"CD",X"D0",X"A4",
		X"C9",X"CD",X"C0",X"3E",X"21",X"16",X"4E",X"CD",X"60",X"8C",X"CD",X"86",X"8C",X"3E",X"03",X"32",
		X"80",X"50",X"CD",X"DB",X"80",X"CD",X"EE",X"80",X"C9",X"3A",X"FE",X"4D",X"A7",X"28",X"07",X"AF",
		X"32",X"FE",X"4D",X"CD",X"B3",X"8D",X"3A",X"FF",X"4D",X"A7",X"C8",X"AF",X"32",X"FF",X"4D",X"CD",
		X"B3",X"8D",X"C9",X"3A",X"A5",X"4D",X"A7",X"C0",X"21",X"FB",X"4D",X"7E",X"A7",X"C8",X"35",X"CD",
		X"49",X"8C",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"C3",X"9C",X"A6",X"78",X"FE",X"05",
		X"20",X"02",X"3D",X"05",X"32",X"A4",X"4D",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3A",X"EA",X"90",X"A7",X"20",X"04",
		X"21",X"3E",X"3D",X"C9",X"21",X"F7",X"8B",X"C9",X"CD",X"A6",X"8E",X"21",X"00",X"90",X"06",X"0F",
		X"AF",X"CF",X"21",X"00",X"00",X"22",X"F0",X"90",X"22",X"F2",X"90",X"C9",X"F5",X"ED",X"57",X"B7",
		X"28",X"04",X"F1",X"C3",X"D4",X"3B",X"F1",X"C3",X"30",X"3D",X"FF",X"CD",X"C2",X"1F",X"3E",X"5C",
		X"32",X"9D",X"41",X"3E",X"01",X"32",X"9D",X"45",X"06",X"17",X"CD",X"5E",X"2C",X"C9",X"FF",X"FF",
		X"FF",X"FF",X"CD",X"51",X"8C",X"3A",X"13",X"4E",X"A7",X"C0",X"CD",X"00",X"81",X"C9",X"FF",X"FF",
		X"06",X"01",X"CD",X"ED",X"23",X"CD",X"D7",X"24",X"CD",X"B3",X"8D",X"AF",X"21",X"E0",X"4D",X"06",
		X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",X"CF",X"CD",X"81",X"8D",X"CD",X"7F",X"0F",X"CD",X"08",
		X"8E",X"CD",X"77",X"25",X"C9",X"06",X"03",X"CD",X"5A",X"2A",X"CD",X"D2",X"8A",X"C3",X"40",X"19",
		X"FE",X"03",X"CA",X"C2",X"8B",X"3E",X"01",X"32",X"E2",X"90",X"C9",X"AF",X"21",X"E0",X"4D",X"06",
		X"20",X"CF",X"21",X"A4",X"4D",X"06",X"0C",X"CF",X"C9",X"FF",X"3E",X"01",X"32",X"80",X"50",X"3A",
		X"F6",X"4D",X"C9",X"CD",X"C0",X"3E",X"3A",X"1C",X"4E",X"CD",X"19",X"81",X"C9",X"3A",X"E4",X"4D",
		X"FE",X"01",X"CA",X"76",X"01",X"FE",X"02",X"28",X"06",X"CD",X"9E",X"84",X"C3",X"76",X"01",X"CD",
		X"D0",X"8E",X"C3",X"76",X"01",X"AF",X"32",X"E4",X"4D",X"CD",X"CC",X"81",X"CD",X"8B",X"87",X"C9",
		X"2A",X"22",X"4C",X"ED",X"5B",X"2A",X"4C",X"22",X"2A",X"4C",X"ED",X"53",X"22",X"4C",X"CD",X"64",
		X"8F",X"ED",X"5B",X"3A",X"4C",X"22",X"3A",X"4C",X"ED",X"53",X"32",X"4C",X"C9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"21",X"48",X"4D",X"7E",X"8F",X"77",X"C9",X"21",X"4C",
		X"3E",X"9E",X"21",X"11",X"42",X"CD",X"DE",X"3C",X"3E",X"01",X"CD",X"F4",X"3C",X"C9",X"FF",X"FF",
		X"CD",X"9E",X"85",X"CD",X"10",X"81",X"C9",X"CD",X"66",X"8D",X"CD",X"A6",X"0A",X"3A",X"09",X"4E",
		X"EE",X"01",X"32",X"09",X"4E",X"C3",X"6C",X"09",X"3A",X"01",X"90",X"A7",X"28",X"07",X"78",X"FE",
		X"04",X"C8",X"FE",X"03",X"C8",X"3A",X"02",X"90",X"A7",X"38",X"07",X"78",X"FE",X"02",X"C8",X"FE",
		X"01",X"C8",X"CD",X"CF",X"88",X"C9",X"3A",X"03",X"90",X"A7",X"28",X"07",X"78",X"FE",X"04",X"C8",
		X"FE",X"03",X"C8",X"3A",X"04",X"90",X"A7",X"28",X"07",X"78",X"FE",X"02",X"C8",X"FE",X"01",X"C8",
		X"CD",X"CF",X"88",X"C9",X"21",X"32",X"4C",X"34",X"2A",X"32",X"4C",X"C9",X"CA",X"B6",X"8B",X"05",
		X"2A",X"D2",X"4D",X"3E",X"10",X"95",X"ED",X"5B",X"08",X"4D",X"A7",X"ED",X"52",X"CA",X"B6",X"8B",
		X"C3",X"08",X"3B",X"3E",X"01",X"32",X"A8",X"4D",X"32",X"AD",X"4D",X"C9",X"CD",X"70",X"84",X"0E",
		X"03",X"3E",X"76",X"21",X"BC",X"41",X"CD",X"DE",X"3C",X"F5",X"3E",X"01",X"CD",X"F4",X"3C",X"F1",
		X"06",X"04",X"80",X"11",X"40",X"00",X"19",X"0D",X"20",X"EC",X"CD",X"2B",X"8E",X"C9",X"00",X"00",
		X"C4",X"40",X"16",X"0F",X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"6C",X"08",X"07",X"00",X"00",X"06",
		X"05",X"00",X"04",X"03",X"02",X"01",X"FE",X"2D",X"2C",X"2B",X"2A",X"29",X"28",X"6D",X"1F",X"1E",
		X"1D",X"1C",X"00",X"00",X"00",X"1B",X"00",X"1A",X"19",X"18",X"17",X"FE",X"6B",X"6A",X"69",X"68",
		X"67",X"66",X"65",X"64",X"63",X"62",X"61",X"00",X"00",X"60",X"3F",X"3E",X"3D",X"3C",X"2F",X"2E",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"4E",X"FE",X"03",X"C0",X"3A",X"04",X"4E",X"FE",X"09",X"28",X"0A",X"FE",X"20",X"20",
		X"06",X"3E",X"01",X"32",X"80",X"50",X"C9",X"3A",X"C1",X"50",X"E6",X"01",X"28",X"30",X"3A",X"E4",
		X"4D",X"A7",X"20",X"1A",X"3A",X"A5",X"4D",X"A7",X"C0",X"3A",X"1C",X"4E",X"A7",X"C8",X"3E",X"01",
		X"32",X"FC",X"90",X"3E",X"70",X"CD",X"9E",X"3E",X"3E",X"05",X"CD",X"AB",X"3E",X"C9",X"FE",X"01",
		X"CA",X"42",X"A1",X"FE",X"02",X"CA",X"D8",X"A3",X"FE",X"03",X"CA",X"83",X"81",X"C9",X"3A",X"FC",
		X"90",X"A7",X"C8",X"AF",X"32",X"FC",X"90",X"3E",X"72",X"CD",X"9E",X"3E",X"3E",X"11",X"CD",X"AB",
		X"3E",X"3A",X"A5",X"4D",X"A7",X"C0",X"3A",X"E4",X"4D",X"A7",X"C8",X"FE",X"03",X"30",X"04",X"CD",
		X"F3",X"A3",X"C9",X"3A",X"F4",X"90",X"A7",X"20",X"03",X"CD",X"AC",X"82",X"AF",X"32",X"E4",X"4D",
		X"32",X"E6",X"4D",X"32",X"F4",X"90",X"32",X"FA",X"4D",X"CD",X"8B",X"87",X"CD",X"5E",X"81",X"C9",
		X"DD",X"21",X"00",X"4C",X"FD",X"21",X"61",X"3E",X"21",X"A7",X"4D",X"06",X"04",X"0E",X"01",X"7E",
		X"A7",X"E5",X"28",X"2B",X"21",X"EF",X"90",X"59",X"16",X"00",X"19",X"7E",X"FE",X"F0",X"28",X"1F",
		X"79",X"87",X"5F",X"DD",X"E5",X"FD",X"E5",X"FD",X"19",X"DD",X"19",X"FD",X"5E",X"00",X"FD",X"23",
		X"FD",X"56",X"00",X"DD",X"73",X"00",X"DD",X"23",X"DD",X"72",X"00",X"FD",X"E1",X"DD",X"E1",X"E1",
		X"23",X"0C",X"05",X"20",X"CA",X"C9",X"3A",X"00",X"4E",X"FE",X"01",X"C8",X"3A",X"04",X"4E",X"FE",
		X"10",X"D0",X"3A",X"72",X"4E",X"4F",X"3A",X"09",X"4E",X"A1",X"28",X"0C",X"3A",X"40",X"50",X"CB",
		X"67",X"28",X"11",X"CD",X"FB",X"A3",X"C9",X"FF",X"3A",X"00",X"50",X"CB",X"77",X"28",X"05",X"CD",
		X"FB",X"A3",X"C9",X"FF",X"3A",X"FB",X"90",X"A7",X"C0",X"3E",X"01",X"32",X"FB",X"90",X"2A",X"EB",
		X"4D",X"3E",X"40",X"77",X"2A",X"39",X"4D",X"CD",X"65",X"00",X"CD",X"58",X"8D",X"22",X"EB",X"4D",
		X"2A",X"39",X"4D",X"22",X"E9",X"4D",X"3A",X"F5",X"90",X"A7",X"C0",X"21",X"BC",X"4E",X"36",X"80",
		X"3E",X"01",X"32",X"F5",X"90",X"C9",X"3A",X"13",X"4E",X"A7",X"C8",X"3A",X"ED",X"90",X"C3",X"DE",
		X"A3",X"FF",X"21",X"9C",X"4E",X"36",X"04",X"CD",X"99",X"8D",X"2A",X"08",X"4D",X"CD",X"83",X"31",
		X"C9",X"21",X"9C",X"4E",X"36",X"08",X"CD",X"99",X"8D",X"2A",X"00",X"4D",X"CD",X"83",X"31",X"C9",
		X"40",X"20",X"CC",X"86",X"77",X"1C",X"0F",X"FF",X"70",X"00",X"01",X"0F",X"00",X"01",X"0C",X"00",
		X"70",X"00",X"01",X"0C",X"00",X"01",X"0C",X"00",X"60",X"00",X"01",X"0C",X"00",X"01",X"0C",X"00",
		X"40",X"00",X"87",X"17",X"00",X"01",X"0C",X"00",X"60",X"A0",X"CC",X"10",X"10",X"02",X"04",X"00",
		X"70",X"20",X"FF",X"86",X"FE",X"1C",X"0F",X"EE",X"31",X"10",X"01",X"0C",X"00",X"01",X"0C",X"00",
		X"3A",X"00",X"4E",X"E7",X"AC",X"A1",X"80",X"A2",X"00",X"A2",X"0E",X"A2",X"3A",X"01",X"4E",X"E7",
		X"5E",X"A2",X"0C",X"00",X"3A",X"02",X"4E",X"E7",X"5D",X"85",X"0C",X"00",X"95",X"A2",X"0C",X"00",
		X"9E",X"A2",X"0C",X"00",X"A7",X"A2",X"0C",X"00",X"AE",X"A2",X"0C",X"00",X"B4",X"A2",X"0C",X"00",
		X"BD",X"A2",X"0C",X"00",X"C4",X"A2",X"0C",X"00",X"CA",X"A2",X"0C",X"00",X"D0",X"A2",X"0C",X"00",
		X"D9",X"A2",X"0C",X"00",X"E0",X"A2",X"0C",X"00",X"E6",X"A2",X"0C",X"00",X"44",X"82",X"0C",X"00",
		X"EF",X"A2",X"0C",X"00",X"F5",X"A2",X"0C",X"00",X"07",X"05",X"0C",X"00",X"EA",X"04",X"7C",X"05",
		X"3A",X"03",X"4E",X"E7",X"0F",X"A3",X"04",X"0A",X"2B",X"32",X"8F",X"06",X"AC",X"06",X"3A",X"04",
		X"4E",X"E7",X"79",X"08",X"99",X"08",X"CD",X"08",X"CD",X"08",X"0D",X"09",X"0C",X"00",X"40",X"09",
		X"0C",X"00",X"EE",X"31",X"A0",X"03",X"0C",X"00",X"D2",X"09",X"D8",X"09",X"0C",X"00",X"E8",X"09",
		X"0C",X"00",X"0B",X"0A",X"0C",X"00",X"02",X"0A",X"0C",X"00",X"04",X"0A",X"0C",X"00",X"06",X"0A",
		X"0C",X"00",X"08",X"0A",X"0C",X"00",X"0A",X"0A",X"0C",X"00",X"0C",X"0A",X"0C",X"00",X"0E",X"0A",
		X"0C",X"00",X"2C",X"0A",X"0C",X"00",X"7C",X"0A",X"A0",X"0A",X"0C",X"00",X"A3",X"0A",X"EF",X"00",
		X"00",X"EF",X"06",X"00",X"EF",X"01",X"00",X"EF",X"14",X"00",X"EF",X"18",X"00",X"EF",X"04",X"00",
		X"EF",X"1E",X"00",X"EF",X"07",X"00",X"21",X"01",X"4E",X"34",X"21",X"C0",X"50",X"36",X"01",X"C9",
		X"CD",X"A1",X"2B",X"3A",X"6E",X"4E",X"A7",X"C3",X"BA",X"A3",X"32",X"04",X"4E",X"32",X"02",X"4E",
		X"21",X"00",X"4E",X"34",X"C9",X"06",X"02",X"CD",X"5E",X"2C",X"CD",X"8A",X"05",X"C9",X"06",X"0C",
		X"CD",X"5E",X"2C",X"CD",X"8A",X"05",X"C9",X"CD",X"D7",X"84",X"CD",X"8A",X"05",X"C9",X"06",X"0D",
		X"CD",X"97",X"A2",X"C9",X"06",X"0E",X"CD",X"97",X"A2",X"CD",X"3E",X"85",X"C9",X"CD",X"ED",X"84",
		X"CD",X"8A",X"05",X"C9",X"06",X"0F",X"CD",X"97",X"A2",X"C9",X"06",X"10",X"CD",X"97",X"A2",X"C9",
		X"06",X"11",X"CD",X"97",X"A2",X"CD",X"45",X"85",X"C9",X"CD",X"F7",X"84",X"CD",X"8A",X"05",X"C9",
		X"06",X"12",X"CD",X"97",X"A2",X"C9",X"06",X"13",X"CD",X"97",X"A2",X"CD",X"4C",X"85",X"C9",X"06",
		X"14",X"CD",X"97",X"A2",X"C9",X"06",X"15",X"CD",X"97",X"A2",X"CD",X"53",X"85",X"C9",X"C9",X"06",
		X"15",X"CD",X"97",X"A2",X"C9",X"80",X"05",X"EF",X"1C",X"11",X"0E",X"12",X"C3",X"85",X"05",X"CD",
		X"A1",X"2B",X"EF",X"00",X"01",X"EF",X"01",X"00",X"EF",X"1C",X"07",X"EF",X"1C",X"0B",X"EF",X"1E",
		X"00",X"21",X"03",X"4E",X"34",X"3E",X"01",X"32",X"D6",X"4D",X"3A",X"71",X"4E",X"FE",X"FF",X"C8",
		X"EF",X"1C",X"0A",X"EF",X"1F",X"00",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"47",X"87",
		X"87",X"80",X"80",X"5F",X"16",X"00",X"DD",X"19",X"DD",X"7E",X"00",X"87",X"47",X"87",X"87",X"4F",
		X"87",X"87",X"81",X"80",X"5F",X"16",X"00",X"21",X"0F",X"33",X"19",X"CD",X"14",X"08",X"DD",X"7E",
		X"01",X"32",X"B0",X"4D",X"DD",X"7E",X"02",X"47",X"87",X"80",X"5F",X"16",X"00",X"21",X"43",X"08",
		X"19",X"CD",X"3A",X"08",X"DD",X"7E",X"03",X"87",X"5F",X"16",X"00",X"FD",X"21",X"4F",X"08",X"FD",
		X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"BB",X"4D",X"DD",X"7E",X"04",X"87",X"5F",X"16",
		X"00",X"FD",X"21",X"61",X"08",X"FD",X"19",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"22",X"BD",X"4D",
		X"DD",X"7E",X"05",X"87",X"5F",X"16",X"00",X"FD",X"21",X"73",X"08",X"FD",X"19",X"FD",X"6E",X"00",
		X"FD",X"66",X"01",X"22",X"95",X"4D",X"CD",X"EA",X"2B",X"C9",X"CA",X"B4",X"A1",X"C3",X"89",X"A2",
		X"FF",X"3A",X"EE",X"90",X"A7",X"20",X"0D",X"3E",X"01",X"32",X"EE",X"90",X"3E",X"00",X"32",X"F2",
		X"45",X"32",X"D2",X"45",X"CD",X"D2",X"2F",X"C9",X"CD",X"51",X"A1",X"C3",X"36",X"A1",X"A7",X"C0",
		X"3E",X"01",X"32",X"ED",X"90",X"21",X"DD",X"DD",X"11",X"DD",X"DD",X"22",X"56",X"4D",X"ED",X"53",
		X"58",X"4D",X"C9",X"CD",X"50",X"8E",X"AF",X"32",X"ED",X"90",X"C9",X"3A",X"FB",X"90",X"A7",X"C8",
		X"21",X"EC",X"90",X"7E",X"FE",X"30",X"28",X"02",X"34",X"C9",X"AF",X"32",X"EC",X"90",X"32",X"FB",
		X"90",X"2A",X"EB",X"4D",X"3E",X"40",X"77",X"21",X"00",X"00",X"22",X"E9",X"4D",X"C9",X"21",X"15",
		X"4E",X"35",X"21",X"00",X"00",X"22",X"EB",X"90",X"CD",X"7C",X"0E",X"3A",X"09",X"4E",X"A7",X"C8",
		X"AF",X"32",X"E3",X"90",X"C9",X"3A",X"EA",X"90",X"A7",X"3E",X"02",X"20",X"02",X"3E",X"03",X"32",
		X"80",X"50",X"C9",X"3A",X"E9",X"90",X"A7",X"C8",X"3A",X"C0",X"4D",X"21",X"20",X"01",X"A7",X"28",
		X"03",X"21",X"24",X"01",X"22",X"0A",X"4C",X"C9",X"32",X"02",X"4C",X"3A",X"E9",X"90",X"A7",X"C8",
		X"3A",X"E6",X"90",X"A7",X"C0",X"3A",X"0A",X"4C",X"81",X"32",X"0A",X"4C",X"C9",X"3A",X"00",X"4E",
		X"FE",X"01",X"28",X"19",X"3A",X"E2",X"90",X"A7",X"28",X"13",X"CD",X"41",X"32",X"C8",X"AF",X"32",
		X"E2",X"90",X"32",X"E4",X"90",X"CD",X"49",X"32",X"28",X"03",X"CD",X"53",X"32",X"CD",X"88",X"09",
		X"CD",X"F9",X"31",X"AF",X"32",X"E4",X"90",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"79",X"A7",X"20",X"0A",X"3A",X"EA",X"90",X"A7",X"C2",X"19",X"1A",X"C3",X"C5",X"18",X"3A",X"E3",
		X"90",X"A7",X"C2",X"19",X"1A",X"C3",X"BF",X"18",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"CD",X"86",X"8C",X"3A",X"EA",X"90",X"A7",X"C8",X"21",X"61",X"43",X"22",X"1A",X"4E",X"C9",X"FF",
		X"3A",X"EA",X"90",X"A7",X"CA",X"CA",X"8D",X"3A",X"E9",X"90",X"A7",X"20",X"36",X"2A",X"39",X"4D",
		X"11",X"27",X"34",X"CD",X"11",X"29",X"2A",X"39",X"4D",X"11",X"27",X"34",X"A7",X"ED",X"52",X"20",
		X"09",X"00",X"00",X"00",X"00",X"00",X"CD",X"83",X"81",X"C9",X"2A",X"39",X"4D",X"11",X"22",X"38",
		X"CD",X"11",X"29",X"2A",X"39",X"4D",X"11",X"22",X"38",X"A7",X"ED",X"52",X"C0",X"3E",X"01",X"32",
		X"E9",X"90",X"C9",X"3A",X"E8",X"90",X"A7",X"20",X"1E",X"2A",X"39",X"4D",X"11",X"22",X"23",X"CD",
		X"11",X"29",X"2A",X"39",X"4D",X"11",X"22",X"23",X"A7",X"ED",X"52",X"C0",X"3E",X"01",X"32",X"E8",
		X"90",X"C9",X"ED",X"72",X"EC",X"FF",X"FF",X"2A",X"39",X"4D",X"11",X"3A",X"25",X"CD",X"11",X"29",
		X"2A",X"39",X"4D",X"11",X"3A",X"25",X"A7",X"ED",X"52",X"20",X"17",X"3E",X"01",X"32",X"E7",X"90",
		X"3E",X"11",X"21",X"9B",X"44",X"CD",X"74",X"0F",X"01",X"42",X"A5",X"21",X"9B",X"40",X"CD",X"72",
		X"81",X"C9",X"3A",X"E7",X"90",X"A7",X"C8",X"2A",X"39",X"4D",X"11",X"3E",X"23",X"CD",X"11",X"29",
		X"2A",X"39",X"4D",X"11",X"3E",X"23",X"A7",X"ED",X"52",X"C0",X"3E",X"17",X"21",X"9B",X"44",X"CD",
		X"74",X"0F",X"3E",X"DE",X"21",X"9B",X"40",X"CD",X"74",X"0F",X"01",X"0B",X"00",X"21",X"3E",X"3D",
		X"11",X"16",X"4E",X"ED",X"B0",X"21",X"16",X"4E",X"CD",X"60",X"8C",X"3E",X"01",X"32",X"E6",X"90",
		X"C9",X"F1",X"00",X"F2",X"02",X"F3",X"0A",X"F4",X"00",X"CD",X"F4",X"00",X"8C",X"F4",X"00",X"8D",
		X"F4",X"00",X"8F",X"F4",X"00",X"8D",X"F4",X"00",X"8C",X"F4",X"00",X"8A",X"F4",X"00",X"AD",X"F4",
		X"00",X"8D",X"F4",X"00",X"8A",X"F4",X"00",X"AD",X"F4",X"00",X"AD",X"F4",X"00",X"8C",X"F4",X"00",
		X"8D",X"F4",X"00",X"8A",X"F4",X"00",X"88",X"F4",X"00",X"85",X"F4",X"00",X"86",X"F4",X"00",X"C8",
		X"F4",X"00",X"88",X"F4",X"00",X"86",X"F4",X"00",X"85",X"F4",X"00",X"83",X"F4",X"00",X"85",X"F4",
		X"00",X"86",X"F4",X"00",X"88",X"F4",X"00",X"8A",X"F4",X"00",X"C8",X"F4",X"00",X"88",X"F4",X"00",
		X"8A",X"F4",X"00",X"8C",X"F4",X"00",X"8A",X"F4",X"00",X"88",X"F4",X"00",X"86",X"F4",X"00",X"85",
		X"F4",X"00",X"83",X"F4",X"00",X"85",X"F4",X"00",X"83",X"F4",X"00",X"C1",X"F4",X"00",X"A1",X"30",
		X"F4",X"00",X"81",X"F4",X"00",X"83",X"F4",X"00",X"A5",X"F4",X"00",X"A6",X"F4",X"00",X"C3",X"F4",
		X"00",X"C8",X"F4",X"00",X"A8",X"F4",X"00",X"88",X"70",X"FF",X"F1",X"01",X"F2",X"03",X"F3",X"06",
		X"F4",X"04",X"81",X"70",X"70",X"00",X"F3",X"03",X"F4",X"04",X"41",X"50",X"30",X"F4",X"04",X"41",
		X"50",X"30",X"F4",X"04",X"41",X"50",X"30",X"F3",X"06",X"F4",X"04",X"81",X"70",X"70",X"00",X"F3",
		X"03",X"F4",X"04",X"41",X"50",X"30",X"F4",X"04",X"41",X"50",X"30",X"F4",X"04",X"41",X"50",X"30",
		X"F3",X"06",X"F4",X"04",X"81",X"70",X"70",X"00",X"F3",X"06",X"F4",X"04",X"81",X"70",X"70",X"00",
		X"F3",X"06",X"F4",X"04",X"81",X"70",X"70",X"00",X"F0",X"56",X"A6",X"FF",X"3A",X"A5",X"4D",X"A7",
		X"28",X"08",X"AF",X"32",X"E5",X"4D",X"32",X"E1",X"90",X"C9",X"3A",X"E5",X"4D",X"A7",X"20",X"19",
		X"2A",X"39",X"4D",X"11",X"3A",X"3A",X"CD",X"11",X"29",X"2A",X"39",X"4D",X"11",X"3A",X"3A",X"A7",
		X"ED",X"52",X"C0",X"3E",X"01",X"32",X"E5",X"4D",X"C9",X"2A",X"39",X"4D",X"11",X"2C",X"27",X"CD",
		X"11",X"29",X"2A",X"39",X"4D",X"11",X"2C",X"27",X"A7",X"ED",X"52",X"20",X"06",X"3E",X"01",X"32",
		X"E1",X"90",X"C9",X"3A",X"E1",X"90",X"A7",X"C8",X"3A",X"A9",X"4D",X"A7",X"20",X"0B",X"2A",X"39",
		X"4D",X"ED",X"5B",X"0E",X"4D",X"CD",X"11",X"29",X"C9",X"AF",X"32",X"E5",X"4D",X"C9",X"21",X"C2",
		X"50",X"06",X"08",X"AF",X"77",X"2C",X"10",X"FC",X"21",X"00",X"40",X"06",X"04",X"32",X"00",X"50",
		X"32",X"07",X"50",X"3E",X"40",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F1",X"06",X"04",X"32",X"00",
		X"50",X"AF",X"32",X"07",X"50",X"3E",X"0F",X"77",X"2C",X"20",X"FC",X"24",X"10",X"F0",X"ED",X"56",
		X"3E",X"FA",X"00",X"00",X"AF",X"32",X"07",X"50",X"3C",X"32",X"C2",X"50",X"FB",X"76",X"31",X"C0",
		X"4F",X"CD",X"70",X"80",X"AF",X"21",X"C2",X"50",X"01",X"08",X"08",X"CF",X"21",X"00",X"4C",X"06",
		X"BE",X"CF",X"CF",X"CF",X"CF",X"21",X"40",X"50",X"06",X"40",X"CF",X"32",X"00",X"50",X"CD",X"0D",
		X"24",X"32",X"00",X"50",X"06",X"00",X"CD",X"ED",X"23",X"32",X"00",X"50",X"21",X"C0",X"4C",X"22",
		X"80",X"4C",X"22",X"82",X"4C",X"3E",X"FF",X"06",X"40",X"CF",X"3E",X"01",X"32",X"C2",X"50",X"FB",
		X"2A",X"82",X"4C",X"7E",X"A7",X"FA",X"80",X"A7",X"36",X"FF",X"2C",X"46",X"36",X"FF",X"2C",X"20",
		X"02",X"2E",X"C0",X"22",X"82",X"4C",X"21",X"80",X"A7",X"E5",X"E7",X"ED",X"23",X"D7",X"24",X"19",
		X"24",X"48",X"24",X"64",X"25",X"8B",X"26",X"0D",X"24",X"98",X"26",X"30",X"27",X"6C",X"27",X"A9",
		X"27",X"F1",X"27",X"3B",X"28",X"65",X"28",X"8F",X"28",X"B9",X"28",X"30",X"02",X"A2",X"26",X"C9",
		X"24",X"35",X"2A",X"D0",X"26",X"87",X"24",X"E8",X"23",X"E0",X"A4",X"E0",X"2A",X"5A",X"2A",X"6A",
		X"2B",X"EA",X"2B",X"5E",X"2C",X"A1",X"2B",X"75",X"26",X"B2",X"26",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
